VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LAYER LEF58_CORNERSPACING STRING ;
END PROPERTYDEFINITIONS

CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.0005 ;
USEMINSPACING OBS ON ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.0115 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.50
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.10        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.28        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.50        0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.06 ENDOFLINE 0.06 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.014 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.15 ;
  WIDTH 0.10 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA12_PG
    LAYER Metal1 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via1 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA12_PG

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_E DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_E

VIA VIA23_1ST_W DEFAULT 
    LAYER Metal2 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_W

VIA VIA23_PG
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via2 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA23_PG

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_N DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_N

VIA VIA34_1ST_S DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_S

VIA VIA34_PG
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via3 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA34_PG

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C

VIA VIA45_PG
    LAYER Metal4 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
    LAYER Via4 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
END VIA45_PG

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA56_PG
    LAYER Metal5 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
    LAYER Via5 ;
        RECT -0.150000 -0.150000 -0.100000 -0.100000 ;
        RECT -0.150000 0.100000 -0.100000 0.150000 ;
        RECT 0.100000 0.100000 0.150000 0.150000 ;
        RECT 0.100000 -0.150000 0.150000 -0.100000 ;
    LAYER Metal6 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
END VIA56_PG

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA6_0_HV

VIA VIA67_PG
    LAYER Metal6 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via6 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA67_PG

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
END VIA7_0_VH

VIA VIA78_PG
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via7 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal8 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA78_PG

VIA VIA8_0_HV DEFAULT 
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
    LAYER Via8 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal9 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
END VIA8_0_HV

VIA VIA12_2C_W DEFAULT
    LAYER Metal1 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA12_2C_W

VIA VIA12_2C_CH DEFAULT
    LAYER Metal1 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via1 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA12_2C_CH

VIA VIA12_2C_E DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via1 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA12_2C_E

VIA VIA12_2C_S DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA12_2C_S

VIA VIA12_2C_CV DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via1 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA12_2C_CV

VIA VIA12_2C_N DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via1 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA12_2C_N

VIA VIA23_2C_W DEFAULT
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA23_2C_W

VIA VIA23_2C_CH DEFAULT
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via2 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA23_2C_CH

VIA VIA23_2C_E DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via2 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA23_2C_E

VIA VIA23_2C_S DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA23_2C_S

VIA VIA23_2C_CV DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via2 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA23_2C_CV

VIA VIA23_2C_N DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via2 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA23_2C_N

VIA VIA34_2C_W DEFAULT
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA34_2C_W

VIA VIA34_2C_CH DEFAULT
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via3 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA34_2C_CH

VIA VIA34_2C_E DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via3 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA34_2C_E

VIA VIA34_2C_S DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA34_2C_S

VIA VIA34_2C_CV DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via3 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA34_2C_CV

VIA VIA34_2C_N DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via3 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA34_2C_N

VIA VIA45_2C_W DEFAULT
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA45_2C_W

VIA VIA45_2C_CH DEFAULT
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via4 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA45_2C_CH

VIA VIA45_2C_E DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via4 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA45_2C_E

VIA VIA45_2C_S DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA45_2C_S

VIA VIA45_2C_CV DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via4 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA45_2C_CV

VIA VIA45_2C_N DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via4 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA45_2C_N

VIA VIA56_2C_W DEFAULT
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA56_2C_W

VIA VIA56_2C_CH DEFAULT
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via5 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal6 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA56_2C_CH

VIA VIA56_2C_E DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via5 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA56_2C_E

VIA VIA56_2C_S DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA56_2C_S

VIA VIA56_2C_CV DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via5 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA56_2C_CV

VIA VIA56_2C_N DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via5 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA56_2C_N

VIA VIA67_2C_W DEFAULT
    LAYER Metal6 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
END VIA67_2C_W

VIA VIA67_2C_CH DEFAULT
    LAYER Metal6 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
    LAYER Via6 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
END VIA67_2C_CH

VIA VIA67_2C_E DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
    LAYER Via6 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
END VIA67_2C_E

VIA VIA67_2C_S DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
END VIA67_2C_S

VIA VIA67_2C_CV DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
    LAYER Via6 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
END VIA67_2C_CV

VIA VIA67_2C_N DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
    LAYER Via6 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
END VIA67_2C_N

VIA VIA78_2C_W DEFAULT
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
END VIA78_2C_W

VIA VIA78_2C_CH DEFAULT
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
    LAYER Via7 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
END VIA78_2C_CH

VIA VIA78_2C_E DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
    LAYER Via7 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
END VIA78_2C_E

VIA VIA78_2C_S DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
END VIA78_2C_S

VIA VIA78_2C_CV DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
    LAYER Via7 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
END VIA78_2C_CV

VIA VIA78_2C_N DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
    LAYER Via7 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
END VIA78_2C_N

VIARULE M4_M3 GENERATE DEFAULT
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
END M4_M3

VIARULE M5_M4 GENERATE DEFAULT
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
END M5_M4

VIARULE M6_M5 GENERATE DEFAULT
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
END M6_M5

VIARULE M7_M6 GENERATE DEFAULT
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
END M7_M6

VIARULE M8_M7 GENERATE DEFAULT
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
END M8_M7

SITE CoreSite
  CLASS CORE ;
  SIZE 0.1 BY 1.2 ;
END CoreSite

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.010 BY 23.5000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 23.5000 BY 23.5000 ;
END corner

MACRO XOR2XL
  CLASS CORE ;
  FOREIGN XOR2XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.291 0.279 1.352 0.795 ;
      RECT 1.262 0.279 1.291 0.360 ;
      RECT 1.282 0.573 1.291 0.627 ;
      RECT 1.262 0.714 1.291 0.795 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.350 0.570 0.379 0.625 ;
      RECT 0.289 0.570 0.350 0.761 ;
      RECT 0.232 0.706 0.289 0.761 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.501 0.557 0.542 0.638 ;
      RECT 0.440 0.439 0.501 0.638 ;
      RECT 0.407 0.439 0.440 0.496 ;
      RECT 0.232 0.442 0.407 0.496 ;
      RECT 0.223 0.433 0.232 0.496 ;
      RECT 0.162 0.388 0.223 0.496 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 -0.080 1.400 0.080 ;
      RECT 1.114 -0.080 1.204 0.122 ;
      RECT 0.325 -0.080 1.114 0.080 ;
      RECT 0.235 -0.080 0.325 0.122 ;
      RECT 0.000 -0.080 0.235 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 1.120 1.400 1.280 ;
      RECT 1.114 1.078 1.204 1.280 ;
      RECT 0.305 1.120 1.114 1.280 ;
      RECT 0.215 1.078 0.305 1.280 ;
      RECT 0.000 1.120 0.215 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.187 0.414 1.229 0.495 ;
      RECT 1.126 0.194 1.187 0.495 ;
      RECT 0.786 0.194 1.126 0.249 ;
      RECT 0.973 0.858 1.063 0.990 ;
      RECT 0.974 0.304 1.035 0.789 ;
      RECT 0.902 0.304 0.974 0.358 ;
      RECT 0.916 0.702 0.974 0.789 ;
      RECT 0.664 0.858 0.973 0.913 ;
      RECT 0.427 0.974 0.875 1.029 ;
      RECT 0.725 0.194 0.786 0.802 ;
      RECT 0.447 0.150 0.664 0.205 ;
      RECT 0.603 0.311 0.664 0.913 ;
      RECT 0.477 0.311 0.603 0.365 ;
      RECT 0.477 0.745 0.603 0.826 ;
      RECT 0.386 0.150 0.447 0.246 ;
      RECT 0.366 0.902 0.427 1.029 ;
      RECT 0.138 0.192 0.386 0.246 ;
      RECT 0.138 0.902 0.366 0.957 ;
      RECT 0.101 0.192 0.138 0.320 ;
      RECT 0.101 0.810 0.138 0.957 ;
      RECT 0.077 0.192 0.101 0.957 ;
      RECT 0.040 0.265 0.077 0.901 ;
  END
END XOR2XL

MACRO XOR2X4
  CLASS CORE ;
  FOREIGN XOR2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.725 0.336 2.786 1.033 ;
      RECT 2.679 0.336 2.725 0.417 ;
      RECT 2.684 0.700 2.725 1.033 ;
      RECT 2.679 0.726 2.684 0.839 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.295 0.500 0.398 0.581 ;
      RECT 0.234 0.500 0.295 0.627 ;
      RECT 0.147 0.500 0.234 0.581 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.999 0.550 2.060 0.627 ;
      RECT 1.888 0.550 1.999 0.605 ;
      RECT 1.797 0.524 1.888 0.605 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.952 -0.080 3.000 0.080 ;
      RECT 2.861 -0.080 2.952 0.122 ;
      RECT 2.588 -0.080 2.861 0.080 ;
      RECT 2.497 -0.080 2.588 0.122 ;
      RECT 2.187 -0.080 2.497 0.080 ;
      RECT 2.096 -0.080 2.187 0.122 ;
      RECT 0.834 -0.080 2.096 0.080 ;
      RECT 0.743 -0.080 0.834 0.122 ;
      RECT 0.481 -0.080 0.743 0.080 ;
      RECT 0.390 -0.080 0.481 0.228 ;
      RECT 0.139 -0.080 0.390 0.080 ;
      RECT 0.048 -0.080 0.139 0.228 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.952 1.120 3.000 1.280 ;
      RECT 2.861 1.078 2.952 1.280 ;
      RECT 2.588 1.120 2.861 1.280 ;
      RECT 2.497 1.078 2.588 1.280 ;
      RECT 2.203 1.120 2.497 1.280 ;
      RECT 2.112 1.078 2.203 1.280 ;
      RECT 0.834 1.120 2.112 1.280 ;
      RECT 0.743 1.078 0.834 1.280 ;
      RECT 0.481 1.120 0.743 1.280 ;
      RECT 0.390 0.989 0.481 1.280 ;
      RECT 0.139 1.120 0.390 1.280 ;
      RECT 0.048 0.989 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.608 0.526 2.663 0.607 ;
      RECT 2.547 0.206 2.608 0.607 ;
      RECT 1.995 0.206 2.547 0.261 ;
      RECT 2.345 0.336 2.406 0.805 ;
      RECT 2.316 0.336 2.345 0.449 ;
      RECT 2.316 0.724 2.345 0.805 ;
      RECT 1.802 0.394 2.316 0.449 ;
      RECT 2.250 0.555 2.283 0.636 ;
      RECT 2.189 0.555 2.250 0.996 ;
      RECT 1.802 0.942 2.189 0.996 ;
      RECT 1.904 0.206 1.995 0.298 ;
      RECT 1.904 0.781 1.995 0.862 ;
      RECT 1.610 0.206 1.904 0.261 ;
      RECT 1.627 0.795 1.904 0.850 ;
      RECT 1.713 0.319 1.802 0.449 ;
      RECT 1.711 0.905 1.802 0.996 ;
      RECT 1.711 0.319 1.713 0.731 ;
      RECT 1.651 0.394 1.711 0.731 ;
      RECT 0.943 0.942 1.711 0.996 ;
      RECT 1.417 0.676 1.651 0.731 ;
      RECT 1.519 0.795 1.627 0.887 ;
      RECT 1.574 0.206 1.610 0.317 ;
      RECT 1.512 0.206 1.574 0.435 ;
      RECT 1.242 0.832 1.519 0.887 ;
      RECT 1.242 0.380 1.512 0.435 ;
      RECT 1.326 0.206 1.417 0.305 ;
      RECT 1.326 0.676 1.417 0.757 ;
      RECT 0.652 0.206 1.326 0.261 ;
      RECT 1.225 0.380 1.242 0.887 ;
      RECT 1.180 0.346 1.225 0.887 ;
      RECT 1.131 0.346 1.180 0.435 ;
      RECT 1.134 0.798 1.180 0.887 ;
      RECT 1.023 0.513 1.103 0.608 ;
      RECT 1.023 0.338 1.037 0.419 ;
      RECT 1.023 0.714 1.037 0.795 ;
      RECT 0.961 0.338 1.023 0.795 ;
      RECT 0.947 0.338 0.961 0.419 ;
      RECT 0.947 0.714 0.961 0.795 ;
      RECT 0.881 0.850 0.943 0.996 ;
      RECT 0.652 0.850 0.881 0.905 ;
      RECT 0.591 0.206 0.652 0.905 ;
      RECT 0.561 0.338 0.591 0.419 ;
      RECT 0.561 0.724 0.591 0.805 ;
      RECT 0.310 0.338 0.561 0.393 ;
      RECT 0.310 0.750 0.561 0.805 ;
      RECT 0.219 0.338 0.310 0.419 ;
      RECT 0.219 0.724 0.310 0.805 ;
  END
END XOR2X4

MACRO XOR2X2
  CLASS CORE ;
  FOREIGN XOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.685 0.171 1.748 0.998 ;
      RECT 1.655 0.171 1.685 0.395 ;
      RECT 1.655 0.693 1.685 0.998 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.368 0.564 0.461 0.694 ;
      RECT 0.326 0.639 0.368 0.694 ;
      RECT 0.263 0.639 0.326 0.763 ;
      RECT 0.239 0.706 0.263 0.763 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.869 0.499 0.931 0.585 ;
      RECT 0.686 0.530 0.869 0.585 ;
      RECT 0.637 0.530 0.686 0.630 ;
      RECT 0.574 0.454 0.637 0.630 ;
      RECT 0.229 0.454 0.574 0.508 ;
      RECT 0.166 0.454 0.229 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.533 -0.080 1.800 0.080 ;
      RECT 1.440 -0.080 1.533 0.122 ;
      RECT 0.720 -0.080 1.440 0.080 ;
      RECT 0.627 -0.080 0.720 0.122 ;
      RECT 0.305 -0.080 0.627 0.080 ;
      RECT 0.213 -0.080 0.305 0.122 ;
      RECT 0.000 -0.080 0.213 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.530 1.120 1.800 1.280 ;
      RECT 1.437 1.078 1.530 1.280 ;
      RECT 0.698 1.120 1.437 1.280 ;
      RECT 0.605 0.905 0.698 1.280 ;
      RECT 0.305 1.120 0.605 1.280 ;
      RECT 0.213 0.905 0.305 1.280 ;
      RECT 0.000 1.120 0.213 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.583 0.473 1.621 0.558 ;
      RECT 1.520 0.212 1.583 0.558 ;
      RECT 1.182 0.212 1.520 0.267 ;
      RECT 1.376 0.520 1.439 0.994 ;
      RECT 0.895 0.939 1.376 0.994 ;
      RECT 1.245 0.336 1.308 0.802 ;
      RECT 1.120 0.212 1.182 0.838 ;
      RECT 1.015 0.212 1.120 0.293 ;
      RECT 1.091 0.783 1.120 0.838 ;
      RECT 0.998 0.783 1.091 0.864 ;
      RECT 0.994 0.368 1.057 0.708 ;
      RECT 0.946 0.368 0.994 0.423 ;
      RECT 0.895 0.654 0.994 0.708 ;
      RECT 0.911 0.206 0.946 0.423 ;
      RECT 0.884 0.163 0.911 0.423 ;
      RECT 0.832 0.654 0.895 0.994 ;
      RECT 0.818 0.163 0.884 0.261 ;
      RECT 0.802 0.717 0.832 0.940 ;
      RECT 0.513 0.206 0.818 0.261 ;
      RECT 0.717 0.319 0.810 0.400 ;
      RECT 0.502 0.765 0.802 0.820 ;
      RECT 0.142 0.332 0.717 0.387 ;
      RECT 0.420 0.193 0.513 0.274 ;
      RECT 0.439 0.765 0.502 0.905 ;
      RECT 0.409 0.824 0.439 0.905 ;
      RECT 0.104 0.281 0.142 0.387 ;
      RECT 0.104 0.683 0.142 0.764 ;
      RECT 0.104 0.950 0.138 1.031 ;
      RECT 0.041 0.281 0.104 1.031 ;
  END
END XOR2X2

MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.291 0.279 1.352 0.788 ;
      RECT 1.262 0.279 1.291 0.360 ;
      RECT 1.282 0.573 1.291 0.788 ;
      RECT 1.262 0.707 1.282 0.788 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.350 0.570 0.379 0.625 ;
      RECT 0.289 0.570 0.350 0.761 ;
      RECT 0.232 0.706 0.289 0.761 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.501 0.557 0.542 0.638 ;
      RECT 0.440 0.439 0.501 0.638 ;
      RECT 0.407 0.439 0.440 0.496 ;
      RECT 0.232 0.442 0.407 0.496 ;
      RECT 0.223 0.433 0.232 0.496 ;
      RECT 0.162 0.388 0.223 0.496 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 -0.080 1.400 0.080 ;
      RECT 1.114 -0.080 1.204 0.122 ;
      RECT 0.325 -0.080 1.114 0.080 ;
      RECT 0.235 -0.080 0.325 0.122 ;
      RECT 0.000 -0.080 0.235 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 1.120 1.400 1.280 ;
      RECT 1.114 1.078 1.204 1.280 ;
      RECT 0.305 1.120 1.114 1.280 ;
      RECT 0.215 1.078 0.305 1.280 ;
      RECT 0.000 1.120 0.215 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.187 0.426 1.229 0.507 ;
      RECT 1.126 0.194 1.187 0.507 ;
      RECT 0.797 0.194 1.126 0.249 ;
      RECT 0.973 0.858 1.063 0.974 ;
      RECT 0.974 0.304 1.035 0.789 ;
      RECT 0.912 0.304 0.974 0.358 ;
      RECT 0.927 0.702 0.974 0.789 ;
      RECT 0.664 0.858 0.973 0.913 ;
      RECT 0.427 0.974 0.875 1.029 ;
      RECT 0.736 0.194 0.797 0.802 ;
      RECT 0.447 0.150 0.675 0.205 ;
      RECT 0.603 0.311 0.664 0.913 ;
      RECT 0.477 0.311 0.603 0.365 ;
      RECT 0.477 0.745 0.603 0.826 ;
      RECT 0.386 0.150 0.447 0.246 ;
      RECT 0.366 0.902 0.427 1.029 ;
      RECT 0.138 0.192 0.386 0.246 ;
      RECT 0.138 0.902 0.366 0.957 ;
      RECT 0.101 0.192 0.138 0.313 ;
      RECT 0.101 0.810 0.138 0.957 ;
      RECT 0.077 0.192 0.101 0.957 ;
      RECT 0.040 0.258 0.077 0.901 ;
  END
END XOR2X1

MACRO XNOR2X4
  CLASS CORE ;
  FOREIGN XNOR2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.725 0.336 2.786 1.033 ;
      RECT 2.679 0.336 2.725 0.417 ;
      RECT 2.684 0.700 2.725 1.033 ;
      RECT 2.679 0.726 2.684 0.807 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.295 0.500 0.398 0.581 ;
      RECT 0.234 0.500 0.295 0.627 ;
      RECT 0.147 0.500 0.234 0.581 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.857 0.517 0.947 0.598 ;
      RECT 0.763 0.517 0.857 0.627 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.952 -0.080 3.000 0.080 ;
      RECT 2.861 -0.080 2.952 0.122 ;
      RECT 2.588 -0.080 2.861 0.080 ;
      RECT 2.497 -0.080 2.588 0.122 ;
      RECT 2.187 -0.080 2.497 0.080 ;
      RECT 2.096 -0.080 2.187 0.122 ;
      RECT 0.834 -0.080 2.096 0.080 ;
      RECT 0.743 -0.080 0.834 0.122 ;
      RECT 0.481 -0.080 0.743 0.080 ;
      RECT 0.390 -0.080 0.481 0.228 ;
      RECT 0.139 -0.080 0.390 0.080 ;
      RECT 0.048 -0.080 0.139 0.228 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.952 1.120 3.000 1.280 ;
      RECT 2.861 1.078 2.952 1.280 ;
      RECT 2.588 1.120 2.861 1.280 ;
      RECT 2.497 1.078 2.588 1.280 ;
      RECT 2.203 1.120 2.497 1.280 ;
      RECT 2.112 1.078 2.203 1.280 ;
      RECT 0.834 1.120 2.112 1.280 ;
      RECT 0.743 1.078 0.834 1.280 ;
      RECT 0.481 1.120 0.743 1.280 ;
      RECT 0.390 0.989 0.481 1.280 ;
      RECT 0.139 1.120 0.390 1.280 ;
      RECT 0.048 0.989 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.608 0.526 2.663 0.607 ;
      RECT 2.547 0.206 2.608 0.961 ;
      RECT 1.995 0.206 2.547 0.261 ;
      RECT 1.134 0.906 2.547 0.961 ;
      RECT 2.345 0.336 2.406 0.805 ;
      RECT 2.316 0.336 2.345 0.449 ;
      RECT 2.316 0.724 2.345 0.805 ;
      RECT 2.037 0.394 2.316 0.449 ;
      RECT 2.250 0.555 2.283 0.636 ;
      RECT 2.189 0.555 2.250 0.851 ;
      RECT 0.652 0.796 2.189 0.851 ;
      RECT 1.976 0.394 2.037 0.715 ;
      RECT 1.904 0.206 1.995 0.298 ;
      RECT 1.802 0.394 1.976 0.449 ;
      RECT 1.417 0.661 1.976 0.715 ;
      RECT 1.610 0.206 1.904 0.261 ;
      RECT 1.797 0.524 1.888 0.605 ;
      RECT 1.723 0.319 1.802 0.449 ;
      RECT 1.070 0.537 1.797 0.592 ;
      RECT 1.711 0.319 1.723 0.400 ;
      RECT 1.574 0.206 1.610 0.317 ;
      RECT 1.512 0.206 1.574 0.401 ;
      RECT 1.134 0.346 1.512 0.401 ;
      RECT 1.326 0.206 1.417 0.292 ;
      RECT 1.326 0.661 1.417 0.742 ;
      RECT 0.652 0.206 1.326 0.261 ;
      RECT 1.008 0.338 1.070 0.733 ;
      RECT 0.947 0.338 1.008 0.419 ;
      RECT 0.947 0.652 1.008 0.733 ;
      RECT 0.591 0.206 0.652 0.851 ;
      RECT 0.561 0.338 0.591 0.419 ;
      RECT 0.561 0.724 0.591 0.805 ;
      RECT 0.310 0.338 0.561 0.393 ;
      RECT 0.310 0.750 0.561 0.805 ;
      RECT 0.219 0.338 0.310 0.419 ;
      RECT 0.219 0.724 0.310 0.805 ;
  END
END XNOR2X4

MACRO XNOR2X2
  CLASS CORE ;
  FOREIGN XNOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.948 0.171 1.950 0.395 ;
      RECT 1.884 0.171 1.948 0.998 ;
      RECT 1.857 0.171 1.884 0.395 ;
      RECT 1.854 0.693 1.884 0.998 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.490 0.564 0.521 0.645 ;
      RECT 0.427 0.564 0.490 0.694 ;
      RECT 0.402 0.627 0.427 0.694 ;
      RECT 0.329 0.639 0.402 0.694 ;
      RECT 0.266 0.639 0.329 0.763 ;
      RECT 0.241 0.706 0.266 0.763 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.059 0.468 1.123 0.585 ;
      RECT 0.875 0.530 1.059 0.585 ;
      RECT 0.811 0.530 0.875 0.630 ;
      RECT 0.668 0.575 0.811 0.630 ;
      RECT 0.647 0.573 0.668 0.630 ;
      RECT 0.584 0.454 0.647 0.630 ;
      RECT 0.231 0.454 0.584 0.508 ;
      RECT 0.168 0.454 0.231 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.741 -0.080 2.000 0.080 ;
      RECT 1.647 -0.080 1.741 0.122 ;
      RECT 0.810 -0.080 1.647 0.080 ;
      RECT 0.716 -0.080 0.810 0.122 ;
      RECT 0.386 -0.080 0.716 0.080 ;
      RECT 0.292 -0.080 0.386 0.122 ;
      RECT 0.000 -0.080 0.292 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.727 1.120 2.000 1.280 ;
      RECT 1.634 1.078 1.727 1.280 ;
      RECT 0.788 1.120 1.634 1.280 ;
      RECT 0.694 0.905 0.788 1.280 ;
      RECT 0.380 1.120 0.694 1.280 ;
      RECT 0.287 0.905 0.380 1.280 ;
      RECT 0.000 1.120 0.287 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.781 0.471 1.820 0.558 ;
      RECT 1.718 0.196 1.781 0.558 ;
      RECT 1.376 0.196 1.718 0.251 ;
      RECT 1.572 0.520 1.635 0.994 ;
      RECT 1.022 0.939 1.572 0.994 ;
      RECT 1.439 0.306 1.503 0.802 ;
      RECT 1.313 0.196 1.376 0.838 ;
      RECT 1.207 0.196 1.313 0.302 ;
      RECT 1.284 0.783 1.313 0.838 ;
      RECT 1.190 0.783 1.284 0.864 ;
      RECT 1.186 0.357 1.249 0.708 ;
      RECT 1.087 0.357 1.186 0.412 ;
      RECT 1.022 0.654 1.186 0.708 ;
      RECT 1.023 0.199 1.087 0.412 ;
      RECT 0.601 0.199 1.023 0.254 ;
      RECT 0.959 0.654 1.022 0.994 ;
      RECT 0.927 0.717 0.959 0.940 ;
      RECT 0.862 0.308 0.956 0.389 ;
      RECT 0.590 0.765 0.927 0.820 ;
      RECT 0.143 0.321 0.862 0.376 ;
      RECT 0.507 0.186 0.601 0.267 ;
      RECT 0.526 0.765 0.590 0.905 ;
      RECT 0.496 0.824 0.526 0.905 ;
      RECT 0.105 0.281 0.143 0.376 ;
      RECT 0.105 0.683 0.143 0.764 ;
      RECT 0.105 0.950 0.139 1.031 ;
      RECT 0.041 0.281 0.105 1.031 ;
  END
END XNOR2X2

MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.291 0.279 1.352 0.788 ;
      RECT 1.262 0.279 1.291 0.360 ;
      RECT 1.282 0.573 1.291 0.788 ;
      RECT 1.262 0.707 1.282 0.788 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.350 0.555 0.379 0.636 ;
      RECT 0.289 0.555 0.350 0.761 ;
      RECT 0.232 0.706 0.289 0.761 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.501 0.557 0.542 0.638 ;
      RECT 0.440 0.439 0.501 0.638 ;
      RECT 0.407 0.439 0.440 0.496 ;
      RECT 0.232 0.442 0.407 0.496 ;
      RECT 0.223 0.439 0.232 0.496 ;
      RECT 0.162 0.388 0.223 0.496 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 -0.080 1.400 0.080 ;
      RECT 1.114 -0.080 1.204 0.122 ;
      RECT 0.325 -0.080 1.114 0.080 ;
      RECT 0.235 -0.080 0.325 0.122 ;
      RECT 0.000 -0.080 0.235 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 1.120 1.400 1.280 ;
      RECT 1.114 1.078 1.204 1.280 ;
      RECT 0.318 1.120 1.114 1.280 ;
      RECT 0.228 1.078 0.318 1.280 ;
      RECT 0.000 1.120 0.228 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.201 0.426 1.229 0.507 ;
      RECT 1.140 0.426 1.201 0.831 ;
      RECT 0.786 0.776 1.140 0.831 ;
      RECT 0.973 0.886 1.063 0.974 ;
      RECT 0.974 0.295 1.035 0.720 ;
      RECT 0.927 0.295 0.974 0.376 ;
      RECT 0.912 0.665 0.974 0.720 ;
      RECT 0.664 0.886 0.973 0.940 ;
      RECT 0.774 0.158 0.864 0.239 ;
      RECT 0.725 0.295 0.786 0.831 ;
      RECT 0.447 0.185 0.774 0.239 ;
      RECT 0.516 0.995 0.719 1.050 ;
      RECT 0.603 0.321 0.664 0.940 ;
      RECT 0.567 0.321 0.603 0.376 ;
      RECT 0.477 0.745 0.603 0.826 ;
      RECT 0.477 0.295 0.567 0.376 ;
      RECT 0.455 0.902 0.516 1.050 ;
      RECT 0.138 0.902 0.455 0.957 ;
      RECT 0.386 0.185 0.447 0.246 ;
      RECT 0.138 0.192 0.386 0.246 ;
      RECT 0.101 0.192 0.138 0.326 ;
      RECT 0.101 0.810 0.138 0.957 ;
      RECT 0.077 0.192 0.101 0.957 ;
      RECT 0.040 0.192 0.077 0.901 ;
  END
END XNOR2X1

MACRO SEDFFXL
  CLASS CORE ;
  FOREIGN SEDFFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.731 0.533 0.873 0.633 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.332 0.543 0.466 0.650 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.583 0.379 4.643 0.824 ;
      RECT 4.518 0.379 4.583 0.433 ;
      RECT 4.505 0.743 4.583 0.824 ;
      RECT 4.428 0.321 4.518 0.433 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.300 0.213 4.361 0.892 ;
      RECT 4.234 0.213 4.300 0.268 ;
      RECT 4.295 0.837 4.300 0.892 ;
      RECT 4.234 0.837 4.295 0.900 ;
      RECT 4.174 0.167 4.234 0.268 ;
      RECT 4.204 0.845 4.234 0.900 ;
      RECT 4.143 0.845 4.204 1.006 ;
      RECT 4.084 0.162 4.174 0.268 ;
      RECT 4.114 0.925 4.143 1.006 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.231 0.839 0.291 0.910 ;
      RECT 0.186 0.855 0.231 0.910 ;
      RECT 0.125 0.855 0.186 0.981 ;
      RECT 0.096 0.900 0.125 0.981 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.055 0.524 1.182 0.627 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.450 0.433 2.574 0.542 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.496 -0.080 4.700 0.080 ;
      RECT 4.406 -0.080 4.496 0.122 ;
      RECT 3.954 -0.080 4.406 0.080 ;
      RECT 3.893 -0.080 3.954 0.358 ;
      RECT 3.230 -0.080 3.893 0.080 ;
      RECT 3.140 -0.080 3.230 0.218 ;
      RECT 2.765 -0.080 3.140 0.080 ;
      RECT 2.676 -0.080 2.765 0.192 ;
      RECT 0.857 -0.080 2.676 0.080 ;
      RECT 0.797 -0.080 0.857 0.199 ;
      RECT 0.174 -0.080 0.797 0.080 ;
      RECT 0.084 -0.080 0.174 0.122 ;
      RECT 0.000 -0.080 0.084 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.536 1.120 4.700 1.280 ;
      RECT 4.432 1.078 4.536 1.280 ;
      RECT 4.002 1.113 4.432 1.280 ;
      RECT 3.913 0.825 4.002 1.280 ;
      RECT 3.296 1.120 3.913 1.280 ;
      RECT 3.048 1.078 3.296 1.280 ;
      RECT 2.759 1.120 3.048 1.280 ;
      RECT 2.363 1.078 2.759 1.280 ;
      RECT 0.778 1.120 2.363 1.280 ;
      RECT 0.688 0.963 0.778 1.280 ;
      RECT 0.372 1.120 0.688 1.280 ;
      RECT 0.282 0.986 0.372 1.280 ;
      RECT 0.000 1.120 0.282 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.205 0.361 4.240 0.758 ;
      RECT 4.184 0.361 4.205 0.771 ;
      RECT 4.179 0.348 4.184 0.771 ;
      RECT 4.095 0.348 4.179 0.429 ;
      RECT 4.116 0.687 4.179 0.771 ;
      RECT 3.893 0.687 4.116 0.742 ;
      RECT 3.816 0.500 4.078 0.581 ;
      RECT 3.803 0.674 3.893 0.755 ;
      RECT 3.756 0.163 3.816 0.581 ;
      RECT 3.791 0.700 3.803 0.755 ;
      RECT 3.731 0.700 3.791 0.994 ;
      RECT 3.503 0.163 3.756 0.218 ;
      RECT 3.669 0.526 3.756 0.581 ;
      RECT 1.786 0.939 3.731 0.994 ;
      RECT 3.547 0.299 3.695 0.354 ;
      RECT 3.628 0.526 3.669 0.815 ;
      RECT 3.608 0.526 3.628 0.855 ;
      RECT 3.567 0.761 3.608 0.855 ;
      RECT 3.505 0.299 3.547 0.658 ;
      RECT 3.487 0.299 3.505 0.870 ;
      RECT 3.445 0.604 3.487 0.870 ;
      RECT 2.585 0.815 3.445 0.870 ;
      RECT 3.323 0.337 3.384 0.746 ;
      RECT 3.062 0.337 3.323 0.392 ;
      RECT 3.054 0.692 3.323 0.746 ;
      RECT 3.173 0.545 3.263 0.626 ;
      RECT 2.933 0.558 3.173 0.613 ;
      RECT 2.972 0.161 3.062 0.400 ;
      RECT 2.826 0.161 2.972 0.215 ;
      RECT 2.863 0.558 2.933 0.738 ;
      RECT 2.825 0.305 2.863 0.738 ;
      RECT 2.802 0.305 2.825 0.721 ;
      RECT 2.335 0.667 2.802 0.721 ;
      RECT 2.681 0.313 2.742 0.513 ;
      RECT 2.615 0.313 2.681 0.368 ;
      RECT 2.554 0.161 2.615 0.368 ;
      RECT 2.495 0.776 2.585 0.870 ;
      RECT 2.177 0.161 2.554 0.215 ;
      RECT 2.214 0.815 2.495 0.870 ;
      RECT 2.426 0.298 2.487 0.379 ;
      RECT 2.214 0.324 2.426 0.379 ;
      RECT 2.275 0.511 2.335 0.721 ;
      RECT 2.154 0.324 2.214 0.870 ;
      RECT 2.117 0.161 2.177 0.264 ;
      RECT 1.837 0.449 2.154 0.504 ;
      RECT 2.113 0.815 2.154 0.870 ;
      RECT 2.011 0.210 2.117 0.264 ;
      RECT 2.064 0.676 2.093 0.757 ;
      RECT 2.003 0.567 2.064 0.757 ;
      RECT 1.982 0.210 2.011 0.290 ;
      RECT 1.757 0.567 2.003 0.621 ;
      RECT 1.921 0.210 1.982 0.392 ;
      RECT 1.757 0.337 1.921 0.392 ;
      RECT 1.792 0.676 1.882 0.757 ;
      RECT 1.734 0.227 1.800 0.282 ;
      RECT 1.634 0.702 1.792 0.757 ;
      RECT 1.725 0.833 1.786 0.994 ;
      RECT 1.696 0.337 1.757 0.621 ;
      RECT 1.673 0.163 1.734 0.282 ;
      RECT 1.696 0.833 1.725 0.914 ;
      RECT 1.027 0.163 1.673 0.218 ;
      RECT 1.573 0.702 1.634 1.050 ;
      RECT 1.219 0.995 1.573 1.050 ;
      RECT 1.422 0.835 1.511 0.940 ;
      RECT 1.414 0.413 1.501 0.514 ;
      RECT 0.736 0.298 1.441 0.352 ;
      RECT 0.628 0.835 1.422 0.889 ;
      RECT 1.353 0.413 1.414 0.780 ;
      RECT 0.613 0.413 1.353 0.468 ;
      RECT 1.299 0.725 1.353 0.780 ;
      RECT 1.158 0.956 1.219 1.050 ;
      RECT 1.047 0.956 1.158 1.011 ;
      RECT 0.940 0.695 1.030 0.776 ;
      RECT 0.636 0.708 0.940 0.763 ;
      RECT 0.675 0.150 0.736 0.352 ;
      RECT 0.456 0.150 0.675 0.205 ;
      RECT 0.546 0.550 0.636 0.763 ;
      RECT 0.567 0.835 0.628 0.979 ;
      RECT 0.553 0.260 0.613 0.468 ;
      RECT 0.477 0.898 0.567 0.979 ;
      RECT 0.137 0.260 0.553 0.314 ;
      RECT 0.506 0.708 0.546 0.763 ;
      RECT 0.446 0.708 0.506 0.788 ;
      RECT 0.431 0.376 0.492 0.467 ;
      RECT 0.262 0.708 0.446 0.763 ;
      RECT 0.262 0.412 0.431 0.467 ;
      RECT 0.202 0.412 0.262 0.763 ;
      RECT 0.123 0.260 0.137 0.424 ;
      RECT 0.123 0.707 0.137 0.788 ;
      RECT 0.076 0.260 0.123 0.788 ;
      RECT 0.062 0.343 0.076 0.788 ;
      RECT 0.047 0.343 0.062 0.424 ;
      RECT 0.047 0.707 0.062 0.788 ;
  END
END SEDFFXL

MACRO SEDFFX4
  CLASS CORE ;
  FOREIGN SEDFFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.885 0.529 1.042 0.633 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.343 0.543 0.524 0.627 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.714 0.332 5.866 0.413 ;
      RECT 5.709 0.690 5.823 0.771 ;
      RECT 5.709 0.300 5.714 0.633 ;
      RECT 5.619 0.300 5.709 0.771 ;
      RECT 5.614 0.300 5.619 0.633 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.535 0.300 5.540 0.633 ;
      RECT 5.445 0.300 5.535 0.771 ;
      RECT 5.440 0.300 5.445 0.633 ;
      RECT 5.395 0.690 5.445 0.771 ;
      RECT 5.439 0.331 5.440 0.412 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.265 0.839 0.292 0.894 ;
      RECT 0.205 0.839 0.265 0.955 ;
      RECT 0.195 0.900 0.205 0.955 ;
      RECT 0.106 0.900 0.195 0.981 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.307 0.573 1.338 0.627 ;
      RECT 1.203 0.573 1.307 0.694 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.572 0.433 2.752 0.529 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.052 -0.080 6.100 0.080 ;
      RECT 5.963 -0.080 6.052 0.247 ;
      RECT 5.697 -0.080 5.963 0.080 ;
      RECT 5.608 -0.080 5.697 0.221 ;
      RECT 5.358 -0.080 5.608 0.080 ;
      RECT 5.268 -0.080 5.358 0.212 ;
      RECT 4.983 -0.080 5.268 0.080 ;
      RECT 4.893 -0.080 4.983 0.385 ;
      RECT 4.255 -0.080 4.893 0.080 ;
      RECT 4.166 -0.080 4.255 0.122 ;
      RECT 3.569 -0.080 4.166 0.080 ;
      RECT 3.479 -0.080 3.569 0.225 ;
      RECT 2.942 -0.080 3.479 0.080 ;
      RECT 2.852 -0.080 2.942 0.223 ;
      RECT 0.902 -0.080 2.852 0.080 ;
      RECT 0.812 -0.080 0.902 0.216 ;
      RECT 0.169 -0.080 0.812 0.080 ;
      RECT 0.079 -0.080 0.169 0.122 ;
      RECT 0.000 -0.080 0.079 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.002 1.120 6.100 1.280 ;
      RECT 5.913 0.965 6.002 1.280 ;
      RECT 5.654 1.120 5.913 1.280 ;
      RECT 5.564 0.989 5.654 1.280 ;
      RECT 5.316 1.120 5.564 1.280 ;
      RECT 5.226 0.989 5.316 1.280 ;
      RECT 4.925 1.120 5.226 1.280 ;
      RECT 4.811 1.078 4.925 1.280 ;
      RECT 4.178 1.120 4.811 1.280 ;
      RECT 4.088 1.078 4.178 1.280 ;
      RECT 3.424 1.120 4.088 1.280 ;
      RECT 3.334 1.078 3.424 1.280 ;
      RECT 2.827 1.120 3.334 1.280 ;
      RECT 2.737 1.078 2.827 1.280 ;
      RECT 2.482 1.120 2.737 1.280 ;
      RECT 2.392 1.078 2.482 1.280 ;
      RECT 0.864 1.120 2.392 1.280 ;
      RECT 0.774 0.941 0.864 1.280 ;
      RECT 0.462 1.120 0.774 1.280 ;
      RECT 0.372 0.920 0.462 1.280 ;
      RECT 0.000 1.120 0.372 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.944 0.524 5.990 0.605 ;
      RECT 5.883 0.524 5.944 0.881 ;
      RECT 5.777 0.524 5.883 0.605 ;
      RECT 5.285 0.826 5.883 0.881 ;
      RECT 5.225 0.342 5.285 0.881 ;
      RECT 5.173 0.342 5.225 0.396 ;
      RECT 5.126 0.807 5.225 0.881 ;
      RECT 5.083 0.204 5.173 0.396 ;
      RECT 4.974 0.807 5.126 0.888 ;
      RECT 4.852 0.471 5.108 0.552 ;
      RECT 4.913 0.640 4.974 0.994 ;
      RECT 3.960 0.939 4.913 0.994 ;
      RECT 4.830 0.471 4.852 0.870 ;
      RECT 4.792 0.251 4.830 0.870 ;
      RECT 4.769 0.251 4.792 0.526 ;
      RECT 3.814 0.815 4.792 0.870 ;
      RECT 4.604 0.251 4.769 0.306 ;
      RECT 4.624 0.392 4.685 0.704 ;
      RECT 4.337 0.649 4.624 0.704 ;
      RECT 4.514 0.225 4.604 0.306 ;
      RECT 3.907 0.225 4.514 0.280 ;
      RECT 4.439 0.385 4.500 0.471 ;
      RECT 3.572 0.385 4.439 0.439 ;
      RECT 4.248 0.504 4.337 0.704 ;
      RECT 3.693 0.649 4.248 0.704 ;
      RECT 3.899 0.939 3.960 1.050 ;
      RECT 3.817 0.199 3.907 0.280 ;
      RECT 3.586 0.995 3.899 1.050 ;
      RECT 3.754 0.815 3.814 0.940 ;
      RECT 3.632 0.649 3.693 0.870 ;
      RECT 2.209 0.815 3.632 0.870 ;
      RECT 3.525 0.954 3.586 1.050 ;
      RECT 3.511 0.318 3.572 0.732 ;
      RECT 2.307 0.954 3.525 1.008 ;
      RECT 3.368 0.318 3.511 0.373 ;
      RECT 3.132 0.677 3.511 0.732 ;
      RECT 3.388 0.505 3.449 0.607 ;
      RECT 3.071 0.505 3.388 0.560 ;
      RECT 3.289 0.286 3.368 0.373 ;
      RECT 3.228 0.163 3.289 0.373 ;
      RECT 3.183 0.163 3.228 0.218 ;
      RECT 3.071 0.288 3.119 0.407 ;
      RECT 3.058 0.288 3.071 0.727 ;
      RECT 3.010 0.352 3.058 0.727 ;
      RECT 2.362 0.673 3.010 0.727 ;
      RECT 2.889 0.313 2.950 0.555 ;
      RECT 2.791 0.313 2.889 0.368 ;
      RECT 2.730 0.150 2.791 0.368 ;
      RECT 2.161 0.150 2.730 0.205 ;
      RECT 2.580 0.290 2.670 0.371 ;
      RECT 2.412 0.317 2.580 0.371 ;
      RECT 2.352 0.317 2.412 0.437 ;
      RECT 2.301 0.540 2.362 0.727 ;
      RECT 2.209 0.382 2.352 0.437 ;
      RECT 2.246 0.954 2.307 1.039 ;
      RECT 1.760 0.985 2.246 1.039 ;
      RECT 2.148 0.382 2.209 0.886 ;
      RECT 2.132 0.150 2.161 0.295 ;
      RECT 1.957 0.382 2.148 0.437 ;
      RECT 2.110 0.831 2.148 0.886 ;
      RECT 2.101 0.150 2.132 0.327 ;
      RECT 2.072 0.214 2.101 0.327 ;
      RECT 2.033 0.618 2.087 0.773 ;
      RECT 1.887 0.273 2.072 0.327 ;
      RECT 2.027 0.537 2.033 0.773 ;
      RECT 1.973 0.537 2.027 0.673 ;
      RECT 1.887 0.537 1.973 0.592 ;
      RECT 1.582 0.163 1.959 0.218 ;
      RECT 1.822 0.738 1.912 0.819 ;
      RECT 1.826 0.273 1.887 0.592 ;
      RECT 1.697 0.764 1.822 0.819 ;
      RECT 1.636 0.764 1.697 1.006 ;
      RECT 1.479 0.423 1.674 0.477 ;
      RECT 1.225 0.951 1.636 1.006 ;
      RECT 0.750 0.287 1.611 0.342 ;
      RECT 1.521 0.163 1.582 0.231 ;
      RECT 1.385 0.835 1.574 0.889 ;
      RECT 1.171 0.176 1.521 0.231 ;
      RECT 1.418 0.411 1.479 0.754 ;
      RECT 0.628 0.411 1.418 0.465 ;
      RECT 1.386 0.699 1.418 0.754 ;
      RECT 1.324 0.815 1.385 0.889 ;
      RECT 0.663 0.815 1.324 0.870 ;
      RECT 1.135 0.925 1.225 1.006 ;
      RECT 0.757 0.688 1.116 0.743 ;
      RECT 0.757 0.520 0.771 0.601 ;
      RECT 0.696 0.520 0.757 0.761 ;
      RECT 0.689 0.165 0.750 0.342 ;
      RECT 0.681 0.520 0.696 0.601 ;
      RECT 0.520 0.706 0.696 0.761 ;
      RECT 0.549 0.165 0.689 0.220 ;
      RECT 0.602 0.815 0.663 0.979 ;
      RECT 0.568 0.275 0.628 0.465 ;
      RECT 0.573 0.898 0.602 0.979 ;
      RECT 0.137 0.275 0.568 0.330 ;
      RECT 0.430 0.706 0.520 0.800 ;
      RECT 0.281 0.385 0.507 0.439 ;
      RECT 0.281 0.706 0.430 0.761 ;
      RECT 0.220 0.385 0.281 0.761 ;
      RECT 0.123 0.275 0.137 0.424 ;
      RECT 0.077 0.275 0.123 0.800 ;
      RECT 0.062 0.343 0.077 0.800 ;
      RECT 0.048 0.343 0.062 0.424 ;
  END
END SEDFFX4

MACRO SEDFFX2
  CLASS CORE ;
  FOREIGN SEDFFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.741 0.533 0.875 0.633 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.373 0.520 0.498 0.642 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.092 0.306 5.153 0.960 ;
      RECT 5.083 0.306 5.092 0.406 ;
      RECT 5.063 0.736 5.092 0.960 ;
      RECT 5.053 0.325 5.083 0.406 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.797 0.325 4.805 0.439 ;
      RECT 4.790 0.306 4.797 0.439 ;
      RECT 4.759 0.306 4.790 0.706 ;
      RECT 4.730 0.306 4.759 0.762 ;
      RECT 4.717 0.325 4.730 0.439 ;
      RECT 4.698 0.605 4.730 0.762 ;
      RECT 4.715 0.325 4.717 0.406 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.243 0.839 0.290 0.894 ;
      RECT 0.197 0.839 0.243 0.955 ;
      RECT 0.183 0.839 0.197 0.981 ;
      RECT 0.108 0.900 0.183 0.981 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.028 0.537 1.177 0.633 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.463 0.433 2.572 0.564 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.974 -0.080 5.200 0.080 ;
      RECT 4.885 -0.080 4.974 0.221 ;
      RECT 4.448 -0.080 4.885 0.080 ;
      RECT 4.358 -0.080 4.448 0.318 ;
      RECT 3.922 -0.080 4.358 0.080 ;
      RECT 4.357 0.267 4.358 0.317 ;
      RECT 3.833 -0.080 3.922 0.237 ;
      RECT 3.228 -0.080 3.833 0.080 ;
      RECT 3.138 -0.080 3.228 0.190 ;
      RECT 2.760 -0.080 3.138 0.080 ;
      RECT 2.671 -0.080 2.760 0.199 ;
      RECT 0.896 -0.080 2.671 0.080 ;
      RECT 0.806 -0.080 0.896 0.179 ;
      RECT 0.168 -0.080 0.806 0.080 ;
      RECT 0.079 -0.080 0.168 0.122 ;
      RECT 0.000 -0.080 0.079 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.964 1.120 5.200 1.280 ;
      RECT 4.874 0.985 4.964 1.280 ;
      RECT 4.390 1.117 4.874 1.280 ;
      RECT 3.996 1.078 4.390 1.280 ;
      RECT 3.271 1.120 3.996 1.280 ;
      RECT 3.003 1.078 3.271 1.280 ;
      RECT 2.656 1.120 3.003 1.280 ;
      RECT 2.320 1.078 2.656 1.280 ;
      RECT 0.776 1.120 2.320 1.280 ;
      RECT 0.687 0.942 0.776 1.280 ;
      RECT 0.393 1.120 0.687 1.280 ;
      RECT 0.303 0.970 0.393 1.280 ;
      RECT 0.000 1.120 0.303 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.981 0.514 5.032 0.642 ;
      RECT 4.972 0.514 4.981 0.915 ;
      RECT 4.920 0.587 4.972 0.915 ;
      RECT 4.589 0.861 4.920 0.915 ;
      RECT 4.589 0.279 4.606 0.687 ;
      RECT 4.546 0.279 4.589 0.944 ;
      RECT 4.529 0.632 4.546 0.944 ;
      RECT 4.500 0.733 4.529 0.944 ;
      RECT 4.390 0.889 4.500 0.944 ;
      RECT 4.396 0.440 4.457 0.527 ;
      RECT 4.269 0.442 4.396 0.527 ;
      RECT 4.329 0.889 4.390 0.960 ;
      RECT 4.268 0.905 4.329 0.960 ;
      RECT 4.209 0.370 4.269 0.717 ;
      RECT 4.178 0.905 4.268 1.008 ;
      RECT 4.075 0.370 4.209 0.425 ;
      RECT 4.164 0.662 4.209 0.717 ;
      RECT 2.260 0.954 4.178 1.008 ;
      RECT 4.075 0.662 4.164 0.743 ;
      RECT 4.059 0.500 4.148 0.581 ;
      RECT 3.985 0.338 4.075 0.425 ;
      RECT 3.870 0.688 4.075 0.743 ;
      RECT 3.704 0.526 4.059 0.581 ;
      RECT 3.704 0.370 3.985 0.425 ;
      RECT 3.809 0.688 3.870 0.838 ;
      RECT 3.639 0.783 3.809 0.838 ;
      RECT 3.644 0.295 3.704 0.425 ;
      RECT 3.644 0.526 3.704 0.658 ;
      RECT 3.574 0.295 3.644 0.350 ;
      RECT 3.542 0.604 3.644 0.658 ;
      RECT 3.549 0.783 3.639 0.864 ;
      RECT 3.485 0.269 3.574 0.350 ;
      RECT 3.249 0.442 3.572 0.496 ;
      RECT 3.452 0.604 3.542 0.688 ;
      RECT 3.427 0.633 3.452 0.688 ;
      RECT 3.367 0.633 3.427 0.874 ;
      RECT 2.524 0.819 3.367 0.874 ;
      RECT 3.188 0.337 3.249 0.764 ;
      RECT 3.070 0.337 3.188 0.392 ;
      RECT 3.029 0.710 3.188 0.764 ;
      RECT 2.871 0.585 3.127 0.639 ;
      RECT 3.041 0.305 3.070 0.392 ;
      RECT 2.995 0.161 3.041 0.392 ;
      RECT 2.981 0.161 2.995 0.386 ;
      RECT 2.846 0.161 2.981 0.215 ;
      RECT 2.810 0.333 2.871 0.732 ;
      RECT 2.754 0.670 2.810 0.732 ;
      RECT 2.257 0.670 2.754 0.725 ;
      RECT 2.675 0.313 2.735 0.550 ;
      RECT 2.611 0.313 2.675 0.368 ;
      RECT 2.550 0.161 2.611 0.368 ;
      RECT 2.226 0.161 2.550 0.215 ;
      RECT 2.420 0.782 2.524 0.874 ;
      RECT 2.416 0.283 2.477 0.379 ;
      RECT 2.136 0.782 2.420 0.837 ;
      RECT 2.403 0.324 2.416 0.379 ;
      RECT 2.343 0.324 2.403 0.444 ;
      RECT 2.136 0.389 2.343 0.444 ;
      RECT 2.199 0.954 2.260 1.050 ;
      RECT 2.197 0.519 2.257 0.725 ;
      RECT 2.165 0.161 2.226 0.263 ;
      RECT 1.762 0.995 2.199 1.050 ;
      RECT 2.003 0.208 2.165 0.263 ;
      RECT 2.076 0.389 2.136 0.912 ;
      RECT 1.803 0.392 2.076 0.446 ;
      RECT 2.037 0.857 2.076 0.912 ;
      RECT 1.954 0.537 2.014 0.781 ;
      RECT 1.974 0.208 2.003 0.300 ;
      RECT 1.913 0.208 1.974 0.336 ;
      RECT 1.681 0.537 1.954 0.592 ;
      RECT 1.681 0.281 1.913 0.336 ;
      RECT 1.750 0.700 1.840 0.781 ;
      RECT 1.040 0.156 1.792 0.211 ;
      RECT 1.702 0.940 1.762 1.050 ;
      RECT 1.614 0.726 1.750 0.781 ;
      RECT 1.620 0.281 1.681 0.592 ;
      RECT 1.553 0.726 1.614 1.046 ;
      RECT 1.169 0.992 1.553 1.046 ;
      RECT 1.396 0.404 1.542 0.458 ;
      RECT 1.395 0.882 1.493 0.937 ;
      RECT 1.405 0.277 1.434 0.332 ;
      RECT 1.345 0.265 1.405 0.332 ;
      RECT 1.335 0.404 1.396 0.762 ;
      RECT 1.334 0.818 1.395 0.937 ;
      RECT 0.746 0.265 1.345 0.320 ;
      RECT 1.250 0.404 1.335 0.458 ;
      RECT 1.295 0.707 1.335 0.762 ;
      RECT 0.626 0.818 1.334 0.873 ;
      RECT 1.190 0.375 1.250 0.458 ;
      RECT 0.625 0.375 1.190 0.430 ;
      RECT 1.108 0.929 1.169 1.046 ;
      RECT 1.044 0.929 1.108 0.983 ;
      RECT 0.625 0.708 1.026 0.763 ;
      RECT 0.685 0.164 0.746 0.320 ;
      RECT 0.494 0.164 0.685 0.219 ;
      RECT 0.625 0.485 0.664 0.539 ;
      RECT 0.576 0.818 0.626 0.952 ;
      RECT 0.565 0.274 0.625 0.430 ;
      RECT 0.565 0.485 0.625 0.763 ;
      RECT 0.566 0.818 0.576 0.979 ;
      RECT 0.487 0.898 0.566 0.979 ;
      RECT 0.137 0.274 0.565 0.329 ;
      RECT 0.494 0.698 0.565 0.763 ;
      RECT 0.303 0.383 0.504 0.438 ;
      RECT 0.404 0.698 0.494 0.779 ;
      RECT 0.303 0.698 0.404 0.752 ;
      RECT 0.243 0.383 0.303 0.752 ;
      RECT 0.122 0.274 0.137 0.424 ;
      RECT 0.076 0.274 0.122 0.800 ;
      RECT 0.062 0.343 0.076 0.800 ;
      RECT 0.047 0.343 0.062 0.424 ;
  END
END SEDFFX2

MACRO SEDFFX1
  CLASS CORE ;
  FOREIGN SEDFFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.731 0.533 0.873 0.633 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.332 0.543 0.466 0.650 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.583 0.379 4.643 0.824 ;
      RECT 4.518 0.379 4.583 0.433 ;
      RECT 4.505 0.743 4.583 0.824 ;
      RECT 4.428 0.320 4.518 0.433 ;
      RECT 4.427 0.333 4.428 0.433 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.300 0.213 4.361 0.892 ;
      RECT 4.234 0.213 4.300 0.268 ;
      RECT 4.295 0.837 4.300 0.892 ;
      RECT 4.234 0.837 4.295 0.900 ;
      RECT 4.084 0.175 4.234 0.268 ;
      RECT 4.204 0.845 4.234 0.900 ;
      RECT 4.143 0.845 4.204 1.006 ;
      RECT 4.114 0.925 4.143 1.006 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.231 0.839 0.291 0.910 ;
      RECT 0.186 0.855 0.231 0.910 ;
      RECT 0.125 0.855 0.186 0.981 ;
      RECT 0.096 0.900 0.125 0.981 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.055 0.524 1.182 0.627 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.450 0.433 2.574 0.542 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.496 -0.080 4.700 0.080 ;
      RECT 4.406 -0.080 4.496 0.122 ;
      RECT 3.954 -0.080 4.406 0.080 ;
      RECT 3.893 -0.080 3.954 0.341 ;
      RECT 3.230 -0.080 3.893 0.080 ;
      RECT 3.140 -0.080 3.230 0.218 ;
      RECT 2.765 -0.080 3.140 0.080 ;
      RECT 2.676 -0.080 2.765 0.192 ;
      RECT 0.857 -0.080 2.676 0.080 ;
      RECT 0.797 -0.080 0.857 0.199 ;
      RECT 0.174 -0.080 0.797 0.080 ;
      RECT 0.084 -0.080 0.174 0.122 ;
      RECT 0.000 -0.080 0.084 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.536 1.120 4.700 1.280 ;
      RECT 4.432 1.078 4.536 1.280 ;
      RECT 4.002 1.113 4.432 1.280 ;
      RECT 3.913 0.846 4.002 1.280 ;
      RECT 3.294 1.120 3.913 1.280 ;
      RECT 3.046 1.078 3.294 1.280 ;
      RECT 2.759 1.120 3.046 1.280 ;
      RECT 2.363 1.078 2.759 1.280 ;
      RECT 0.778 1.120 2.363 1.280 ;
      RECT 0.688 0.963 0.778 1.280 ;
      RECT 0.372 1.120 0.688 1.280 ;
      RECT 0.282 0.986 0.372 1.280 ;
      RECT 0.000 1.120 0.282 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.184 0.361 4.240 0.752 ;
      RECT 4.179 0.348 4.184 0.752 ;
      RECT 4.095 0.348 4.179 0.429 ;
      RECT 4.116 0.671 4.179 0.752 ;
      RECT 3.893 0.689 4.116 0.744 ;
      RECT 3.816 0.500 4.078 0.581 ;
      RECT 3.803 0.676 3.893 0.757 ;
      RECT 3.756 0.163 3.816 0.581 ;
      RECT 3.791 0.702 3.803 0.757 ;
      RECT 3.731 0.702 3.791 0.994 ;
      RECT 3.503 0.163 3.756 0.218 ;
      RECT 3.669 0.526 3.756 0.581 ;
      RECT 1.786 0.939 3.731 0.994 ;
      RECT 3.547 0.299 3.695 0.354 ;
      RECT 3.608 0.526 3.669 0.815 ;
      RECT 3.567 0.729 3.608 0.815 ;
      RECT 3.505 0.299 3.547 0.658 ;
      RECT 3.487 0.299 3.505 0.870 ;
      RECT 3.445 0.604 3.487 0.870 ;
      RECT 2.968 0.815 3.445 0.870 ;
      RECT 3.323 0.337 3.384 0.746 ;
      RECT 3.062 0.337 3.323 0.392 ;
      RECT 3.054 0.692 3.323 0.746 ;
      RECT 3.173 0.545 3.263 0.626 ;
      RECT 2.933 0.558 3.173 0.613 ;
      RECT 2.972 0.161 3.062 0.400 ;
      RECT 2.826 0.161 2.972 0.215 ;
      RECT 2.585 0.806 2.968 0.870 ;
      RECT 2.863 0.558 2.933 0.738 ;
      RECT 2.858 0.305 2.863 0.738 ;
      RECT 2.802 0.305 2.858 0.613 ;
      RECT 2.335 0.683 2.858 0.738 ;
      RECT 2.681 0.313 2.742 0.513 ;
      RECT 2.615 0.313 2.681 0.368 ;
      RECT 2.554 0.161 2.615 0.368 ;
      RECT 2.495 0.793 2.585 0.874 ;
      RECT 2.177 0.161 2.554 0.215 ;
      RECT 2.214 0.815 2.495 0.870 ;
      RECT 2.426 0.298 2.487 0.379 ;
      RECT 2.214 0.324 2.426 0.379 ;
      RECT 2.275 0.511 2.335 0.738 ;
      RECT 2.154 0.324 2.214 0.870 ;
      RECT 2.117 0.161 2.177 0.264 ;
      RECT 1.837 0.449 2.154 0.504 ;
      RECT 2.113 0.815 2.154 0.870 ;
      RECT 2.011 0.210 2.117 0.264 ;
      RECT 2.064 0.676 2.093 0.757 ;
      RECT 2.003 0.567 2.064 0.757 ;
      RECT 1.982 0.210 2.011 0.290 ;
      RECT 1.757 0.567 2.003 0.621 ;
      RECT 1.921 0.210 1.982 0.392 ;
      RECT 1.757 0.337 1.921 0.392 ;
      RECT 1.792 0.676 1.882 0.757 ;
      RECT 1.734 0.227 1.800 0.282 ;
      RECT 1.634 0.702 1.792 0.757 ;
      RECT 1.725 0.833 1.786 0.994 ;
      RECT 1.696 0.337 1.757 0.621 ;
      RECT 1.673 0.163 1.734 0.282 ;
      RECT 1.696 0.833 1.725 0.914 ;
      RECT 1.027 0.163 1.673 0.218 ;
      RECT 1.573 0.702 1.634 1.050 ;
      RECT 1.219 0.995 1.573 1.050 ;
      RECT 1.422 0.835 1.511 0.940 ;
      RECT 1.414 0.413 1.501 0.514 ;
      RECT 0.736 0.298 1.441 0.352 ;
      RECT 0.628 0.835 1.422 0.889 ;
      RECT 1.353 0.413 1.414 0.780 ;
      RECT 0.613 0.413 1.353 0.468 ;
      RECT 1.299 0.725 1.353 0.780 ;
      RECT 1.158 0.956 1.219 1.050 ;
      RECT 1.047 0.956 1.158 1.011 ;
      RECT 0.940 0.695 1.030 0.776 ;
      RECT 0.636 0.708 0.940 0.763 ;
      RECT 0.675 0.150 0.736 0.352 ;
      RECT 0.456 0.150 0.675 0.205 ;
      RECT 0.546 0.550 0.636 0.763 ;
      RECT 0.567 0.835 0.628 0.985 ;
      RECT 0.553 0.260 0.613 0.468 ;
      RECT 0.477 0.921 0.567 1.002 ;
      RECT 0.137 0.260 0.553 0.314 ;
      RECT 0.506 0.708 0.546 0.763 ;
      RECT 0.446 0.708 0.506 0.800 ;
      RECT 0.431 0.376 0.492 0.467 ;
      RECT 0.262 0.708 0.446 0.763 ;
      RECT 0.262 0.412 0.431 0.467 ;
      RECT 0.202 0.412 0.262 0.763 ;
      RECT 0.123 0.260 0.137 0.424 ;
      RECT 0.123 0.719 0.137 0.800 ;
      RECT 0.076 0.260 0.123 0.800 ;
      RECT 0.062 0.343 0.076 0.800 ;
      RECT 0.047 0.343 0.062 0.424 ;
      RECT 0.047 0.719 0.062 0.800 ;
  END
END SEDFFX1

MACRO SEDFFHQX4
  CLASS CORE ;
  FOREIGN SEDFFHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.371 0.167 0.512 0.262 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.170 0.490 0.291 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 6.336 0.433 6.389 0.767 ;
      RECT 6.289 0.345 6.336 0.767 ;
      RECT 6.246 0.345 6.289 0.733 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.774 0.549 1.874 0.693 ;
      RECT 1.704 0.555 1.774 0.610 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.079 0.433 1.180 0.564 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.549 0.494 2.605 0.575 ;
      RECT 2.479 0.494 2.549 0.627 ;
      RECT 2.421 0.494 2.479 0.575 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.514 -0.080 6.600 0.080 ;
      RECT 6.425 -0.080 6.514 0.122 ;
      RECT 6.146 -0.080 6.425 0.080 ;
      RECT 6.057 -0.080 6.146 0.364 ;
      RECT 5.757 -0.080 6.057 0.080 ;
      RECT 5.667 -0.080 5.757 0.122 ;
      RECT 4.425 -0.080 5.667 0.080 ;
      RECT 4.336 -0.080 4.425 0.122 ;
      RECT 4.025 -0.080 4.336 0.080 ;
      RECT 3.936 -0.080 4.025 0.122 ;
      RECT 3.433 -0.080 3.936 0.080 ;
      RECT 3.343 -0.080 3.433 0.287 ;
      RECT 2.733 -0.080 3.343 0.080 ;
      RECT 2.643 -0.080 2.733 0.122 ;
      RECT 1.822 -0.080 2.643 0.080 ;
      RECT 1.733 -0.080 1.822 0.122 ;
      RECT 1.114 -0.080 1.733 0.080 ;
      RECT 1.025 -0.080 1.114 0.122 ;
      RECT 0.295 -0.080 1.025 0.080 ;
      RECT 0.205 -0.080 0.295 0.122 ;
      RECT 0.000 -0.080 0.205 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.517 1.120 6.600 1.280 ;
      RECT 6.428 1.078 6.517 1.280 ;
      RECT 6.146 1.120 6.428 1.280 ;
      RECT 6.057 0.735 6.146 1.280 ;
      RECT 5.757 1.120 6.057 1.280 ;
      RECT 5.530 1.078 5.757 1.280 ;
      RECT 3.220 1.120 5.530 1.280 ;
      RECT 2.978 1.078 3.220 1.280 ;
      RECT 2.701 1.120 2.978 1.280 ;
      RECT 2.612 1.078 2.701 1.280 ;
      RECT 1.818 1.120 2.612 1.280 ;
      RECT 1.729 1.078 1.818 1.280 ;
      RECT 1.112 1.120 1.729 1.280 ;
      RECT 1.022 1.078 1.112 1.280 ;
      RECT 0.311 1.120 1.022 1.280 ;
      RECT 0.221 1.078 0.311 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.938 0.507 6.186 0.589 ;
      RECT 5.938 0.290 5.957 0.371 ;
      RECT 5.942 0.717 5.957 0.910 ;
      RECT 5.938 0.717 5.942 1.007 ;
      RECT 5.878 0.290 5.938 1.007 ;
      RECT 5.867 0.290 5.878 0.371 ;
      RECT 5.867 0.717 5.878 1.007 ;
      RECT 4.338 0.952 5.867 1.007 ;
      RECT 5.747 0.543 5.782 0.627 ;
      RECT 5.687 0.192 5.747 0.898 ;
      RECT 4.920 0.192 5.687 0.246 ;
      RECT 4.793 0.843 5.687 0.898 ;
      RECT 5.563 0.301 5.624 0.787 ;
      RECT 4.784 0.301 5.563 0.356 ;
      RECT 4.983 0.732 5.563 0.787 ;
      RECT 5.430 0.418 5.491 0.586 ;
      RECT 4.732 0.531 5.430 0.586 ;
      RECT 4.571 0.301 4.784 0.392 ;
      RECT 4.671 0.531 4.732 0.898 ;
      RECT 4.551 0.151 4.722 0.206 ;
      RECT 4.625 0.531 4.671 0.586 ;
      RECT 4.211 0.843 4.671 0.898 ;
      RECT 4.550 0.692 4.611 0.787 ;
      RECT 4.211 0.301 4.571 0.356 ;
      RECT 4.491 0.151 4.551 0.246 ;
      RECT 4.211 0.732 4.550 0.787 ;
      RECT 3.821 0.192 4.491 0.246 ;
      RECT 4.278 0.952 4.338 1.050 ;
      RECT 3.363 0.995 4.278 1.050 ;
      RECT 4.150 0.301 4.211 0.787 ;
      RECT 4.150 0.843 4.211 0.940 ;
      RECT 3.486 0.886 4.150 0.940 ;
      RECT 4.013 0.508 4.074 0.831 ;
      RECT 3.608 0.776 4.013 0.831 ;
      RECT 3.745 0.665 3.836 0.720 ;
      RECT 3.745 0.192 3.821 0.355 ;
      RECT 3.684 0.192 3.745 0.720 ;
      RECT 3.547 0.281 3.608 0.831 ;
      RECT 3.311 0.627 3.547 0.682 ;
      RECT 3.426 0.357 3.487 0.549 ;
      RECT 3.425 0.843 3.486 0.940 ;
      RECT 3.093 0.357 3.426 0.412 ;
      RECT 3.147 0.843 3.425 0.898 ;
      RECT 3.303 0.952 3.363 1.050 ;
      RECT 3.250 0.540 3.311 0.682 ;
      RECT 3.025 0.952 3.303 1.007 ;
      RECT 3.087 0.735 3.147 0.898 ;
      RECT 3.033 0.244 3.093 0.680 ;
      RECT 2.909 0.735 3.087 0.789 ;
      RECT 2.986 0.244 3.033 0.299 ;
      RECT 2.986 0.625 3.033 0.680 ;
      RECT 2.964 0.844 3.025 1.007 ;
      RECT 2.909 0.394 2.967 0.449 ;
      RECT 2.329 0.844 2.964 0.899 ;
      RECT 2.849 0.257 2.909 0.789 ;
      RECT 2.453 0.954 2.867 1.008 ;
      RECT 2.528 0.257 2.849 0.312 ;
      RECT 2.412 0.717 2.849 0.771 ;
      RECT 2.438 0.231 2.528 0.312 ;
      RECT 2.392 0.954 2.453 1.031 ;
      RECT 1.967 0.976 2.392 1.031 ;
      RECT 2.316 0.306 2.329 0.899 ;
      RECT 2.268 0.306 2.316 0.915 ;
      RECT 2.226 0.835 2.268 0.915 ;
      RECT 2.161 0.390 2.192 0.742 ;
      RECT 2.139 0.390 2.161 0.888 ;
      RECT 2.132 0.306 2.139 0.888 ;
      RECT 2.079 0.306 2.132 0.445 ;
      RECT 2.126 0.687 2.132 0.888 ;
      RECT 2.100 0.687 2.126 0.915 ;
      RECT 2.037 0.833 2.100 0.915 ;
      RECT 2.018 0.542 2.070 0.631 ;
      RECT 2.018 0.150 2.054 0.205 ;
      RECT 1.437 0.833 2.037 0.888 ;
      RECT 1.958 0.150 2.018 0.749 ;
      RECT 1.907 0.954 1.967 1.031 ;
      RECT 1.613 0.192 1.958 0.246 ;
      RECT 0.670 0.954 1.907 1.008 ;
      RECT 1.832 0.375 1.892 0.482 ;
      RECT 1.613 0.427 1.832 0.482 ;
      RECT 1.613 0.681 1.657 0.736 ;
      RECT 1.613 0.302 1.649 0.357 ;
      RECT 1.553 0.161 1.613 0.246 ;
      RECT 1.553 0.302 1.613 0.736 ;
      RECT 1.299 0.161 1.553 0.215 ;
      RECT 1.521 0.526 1.553 0.613 ;
      RECT 1.376 0.287 1.437 0.888 ;
      RECT 1.008 0.833 1.376 0.888 ;
      RECT 1.242 0.300 1.303 0.725 ;
      RECT 1.172 0.300 1.242 0.355 ;
      RECT 1.172 0.670 1.242 0.725 ;
      RECT 0.947 0.202 1.008 0.888 ;
      RECT 0.889 0.202 0.947 0.257 ;
      RECT 0.797 0.833 0.947 0.888 ;
      RECT 0.829 0.163 0.889 0.257 ;
      RECT 0.825 0.318 0.886 0.733 ;
      RECT 0.797 0.163 0.829 0.218 ;
      RECT 0.786 0.469 0.825 0.554 ;
      RECT 0.670 0.343 0.701 0.501 ;
      RECT 0.641 0.343 0.670 1.008 ;
      RECT 0.609 0.446 0.641 1.008 ;
      RECT 0.470 0.935 0.530 1.050 ;
      RECT 0.476 0.343 0.505 0.424 ;
      RECT 0.476 0.746 0.484 0.827 ;
      RECT 0.416 0.343 0.476 0.827 ;
      RECT 0.137 0.935 0.470 0.989 ;
      RECT 0.395 0.746 0.416 0.827 ;
      RECT 0.108 0.343 0.137 0.424 ;
      RECT 0.108 0.746 0.137 0.989 ;
      RECT 0.076 0.343 0.108 0.989 ;
      RECT 0.047 0.343 0.076 0.827 ;
  END
END SEDFFHQX4

MACRO SEDFFHQX2
  CLASS CORE ;
  FOREIGN SEDFFHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.371 0.167 0.511 0.262 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.170 0.490 0.291 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.862 0.346 5.863 0.733 ;
      RECT 5.803 0.346 5.862 0.767 ;
      RECT 5.758 0.346 5.803 0.427 ;
      RECT 5.763 0.652 5.803 0.767 ;
      RECT 5.758 0.652 5.763 0.733 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.772 0.549 1.872 0.693 ;
      RECT 1.702 0.555 1.772 0.610 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.078 0.433 1.179 0.564 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.448 0.421 2.628 0.512 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.669 -0.080 5.900 0.080 ;
      RECT 5.579 -0.080 5.669 0.122 ;
      RECT 5.294 -0.080 5.579 0.080 ;
      RECT 5.205 -0.080 5.294 0.122 ;
      RECT 4.400 -0.080 5.205 0.080 ;
      RECT 4.311 -0.080 4.400 0.395 ;
      RECT 4.021 -0.080 4.311 0.080 ;
      RECT 3.932 -0.080 4.021 0.342 ;
      RECT 3.430 -0.080 3.932 0.080 ;
      RECT 3.340 -0.080 3.430 0.287 ;
      RECT 2.730 -0.080 3.340 0.080 ;
      RECT 2.641 -0.080 2.730 0.122 ;
      RECT 1.821 -0.080 2.641 0.080 ;
      RECT 1.731 -0.080 1.821 0.122 ;
      RECT 1.113 -0.080 1.731 0.080 ;
      RECT 1.024 -0.080 1.113 0.122 ;
      RECT 0.294 -0.080 1.024 0.080 ;
      RECT 0.205 -0.080 0.294 0.122 ;
      RECT 0.000 -0.080 0.205 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.669 1.120 5.900 1.280 ;
      RECT 5.579 1.078 5.669 1.280 ;
      RECT 5.276 1.120 5.579 1.280 ;
      RECT 5.186 1.078 5.276 1.280 ;
      RECT 3.238 1.120 5.186 1.280 ;
      RECT 3.149 1.078 3.238 1.280 ;
      RECT 2.684 1.120 3.149 1.280 ;
      RECT 2.624 0.902 2.684 1.280 ;
      RECT 1.817 1.120 2.624 1.280 ;
      RECT 1.727 1.078 1.817 1.280 ;
      RECT 1.111 1.120 1.727 1.280 ;
      RECT 1.021 1.078 1.111 1.280 ;
      RECT 0.310 1.120 1.021 1.280 ;
      RECT 0.221 1.078 0.310 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.652 0.500 5.741 0.581 ;
      RECT 5.494 0.526 5.652 0.581 ;
      RECT 5.492 0.292 5.494 0.373 ;
      RECT 5.492 0.526 5.494 0.940 ;
      RECT 5.432 0.292 5.492 0.940 ;
      RECT 5.404 0.292 5.432 0.373 ;
      RECT 5.404 0.748 5.432 0.940 ;
      RECT 5.177 0.855 5.404 0.910 ;
      RECT 5.353 0.543 5.368 0.624 ;
      RECT 5.278 0.543 5.353 0.627 ;
      RECT 5.165 0.573 5.278 0.627 ;
      RECT 5.116 0.683 5.177 0.910 ;
      RECT 5.105 0.213 5.165 0.627 ;
      RECT 5.114 0.855 5.116 0.910 ;
      RECT 5.053 0.855 5.114 1.050 ;
      RECT 5.092 0.213 5.105 0.268 ;
      RECT 5.034 0.573 5.105 0.627 ;
      RECT 5.031 0.174 5.092 0.268 ;
      RECT 3.360 0.995 5.053 1.050 ;
      RECT 4.901 0.330 5.038 0.385 ;
      RECT 4.973 0.573 5.034 0.773 ;
      RECT 4.894 0.174 5.031 0.229 ;
      RECT 4.942 0.718 4.973 0.773 ;
      RECT 4.927 0.718 4.942 0.895 ;
      RECT 4.881 0.718 4.927 0.927 ;
      RECT 4.840 0.330 4.901 0.649 ;
      RECT 4.834 0.150 4.894 0.229 ;
      RECT 4.852 0.814 4.881 0.927 ;
      RECT 4.549 0.873 4.852 0.927 ;
      RECT 4.730 0.594 4.840 0.649 ;
      RECT 4.533 0.150 4.834 0.205 ;
      RECT 4.670 0.737 4.752 0.792 ;
      RECT 4.670 0.261 4.737 0.315 ;
      RECT 4.609 0.261 4.670 0.792 ;
      RECT 4.196 0.470 4.609 0.525 ;
      RECT 4.488 0.735 4.549 0.927 ;
      RECT 4.399 0.594 4.545 0.649 ;
      RECT 4.472 0.150 4.533 0.242 ;
      RECT 4.338 0.594 4.399 0.940 ;
      RECT 3.482 0.886 4.338 0.940 ;
      RECT 4.196 0.276 4.211 0.357 ;
      RECT 4.136 0.276 4.196 0.805 ;
      RECT 4.121 0.276 4.136 0.357 ;
      RECT 4.010 0.508 4.070 0.831 ;
      RECT 3.605 0.776 4.010 0.831 ;
      RECT 3.741 0.289 3.832 0.344 ;
      RECT 3.741 0.665 3.832 0.720 ;
      RECT 3.681 0.289 3.741 0.720 ;
      RECT 3.544 0.231 3.605 0.831 ;
      RECT 3.233 0.554 3.544 0.608 ;
      RECT 3.422 0.843 3.482 0.940 ;
      RECT 3.418 0.357 3.478 0.462 ;
      RECT 2.926 0.843 3.422 0.898 ;
      RECT 3.091 0.357 3.418 0.412 ;
      RECT 3.300 0.954 3.360 1.050 ;
      RECT 2.805 0.954 3.300 1.008 ;
      RECT 3.072 0.268 3.091 0.650 ;
      RECT 3.047 0.255 3.072 0.650 ;
      RECT 3.030 0.255 3.047 0.783 ;
      RECT 2.983 0.255 3.030 0.336 ;
      RECT 2.987 0.595 3.030 0.783 ;
      RECT 2.758 0.394 2.964 0.449 ;
      RECT 2.866 0.665 2.926 0.898 ;
      RECT 2.758 0.665 2.866 0.720 ;
      RECT 2.745 0.776 2.805 1.008 ;
      RECT 2.698 0.257 2.758 0.720 ;
      RECT 2.327 0.776 2.745 0.831 ;
      RECT 2.525 0.257 2.698 0.312 ;
      RECT 2.410 0.665 2.698 0.720 ;
      RECT 2.436 0.231 2.525 0.312 ;
      RECT 1.972 0.982 2.440 1.037 ;
      RECT 2.266 0.306 2.327 0.915 ;
      RECT 2.138 0.390 2.190 0.902 ;
      RECT 2.130 0.306 2.138 0.902 ;
      RECT 2.077 0.306 2.130 0.445 ;
      RECT 2.063 0.833 2.130 0.902 ;
      RECT 2.031 0.542 2.068 0.631 ;
      RECT 1.436 0.833 2.063 0.888 ;
      RECT 2.017 0.150 2.052 0.205 ;
      RECT 2.017 0.542 2.031 0.749 ;
      RECT 1.956 0.150 2.017 0.749 ;
      RECT 1.911 0.954 1.972 1.037 ;
      RECT 1.612 0.192 1.956 0.246 ;
      RECT 1.942 0.668 1.956 0.749 ;
      RECT 0.684 0.954 1.911 1.008 ;
      RECT 1.830 0.375 1.890 0.482 ;
      RECT 1.612 0.427 1.830 0.482 ;
      RECT 1.612 0.668 1.655 0.749 ;
      RECT 1.612 0.302 1.647 0.357 ;
      RECT 1.551 0.161 1.612 0.246 ;
      RECT 1.566 0.302 1.612 0.749 ;
      RECT 1.551 0.302 1.566 0.736 ;
      RECT 1.298 0.161 1.551 0.215 ;
      RECT 1.520 0.526 1.551 0.613 ;
      RECT 1.436 0.287 1.450 0.368 ;
      RECT 1.375 0.287 1.436 0.899 ;
      RECT 1.361 0.287 1.375 0.368 ;
      RECT 1.007 0.844 1.375 0.899 ;
      RECT 1.261 0.300 1.300 0.725 ;
      RECT 1.240 0.287 1.261 0.738 ;
      RECT 1.171 0.287 1.240 0.368 ;
      RECT 1.171 0.657 1.240 0.738 ;
      RECT 0.947 0.202 1.007 0.899 ;
      RECT 0.889 0.202 0.947 0.257 ;
      RECT 0.797 0.844 0.947 0.899 ;
      RECT 0.828 0.163 0.889 0.257 ;
      RECT 0.824 0.318 0.885 0.733 ;
      RECT 0.797 0.163 0.828 0.218 ;
      RECT 0.785 0.469 0.824 0.554 ;
      RECT 0.686 0.343 0.715 0.424 ;
      RECT 0.669 0.343 0.686 0.501 ;
      RECT 0.669 0.820 0.684 1.008 ;
      RECT 0.626 0.343 0.669 1.008 ;
      RECT 0.623 0.446 0.626 1.008 ;
      RECT 0.609 0.446 0.623 0.901 ;
      RECT 0.594 0.820 0.609 0.901 ;
      RECT 0.530 0.969 0.544 1.050 ;
      RECT 0.455 0.935 0.530 1.050 ;
      RECT 0.476 0.343 0.505 0.424 ;
      RECT 0.476 0.746 0.484 0.827 ;
      RECT 0.415 0.343 0.476 0.827 ;
      RECT 0.137 0.935 0.455 0.989 ;
      RECT 0.394 0.746 0.415 0.827 ;
      RECT 0.108 0.343 0.137 0.424 ;
      RECT 0.108 0.746 0.137 0.989 ;
      RECT 0.076 0.343 0.108 0.989 ;
      RECT 0.047 0.343 0.076 0.827 ;
  END
END SEDFFHQX2

MACRO SEDFFHQX1
  CLASS CORE ;
  FOREIGN SEDFFHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.372 0.167 0.513 0.262 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.170 0.490 0.292 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.283 0.324 5.343 0.771 ;
      RECT 5.227 0.324 5.283 0.405 ;
      RECT 5.251 0.690 5.283 0.771 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.779 0.549 1.879 0.693 ;
      RECT 1.709 0.555 1.779 0.610 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.082 0.433 1.184 0.564 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.457 0.421 2.638 0.512 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.169 -0.080 5.400 0.080 ;
      RECT 5.079 -0.080 5.169 0.122 ;
      RECT 4.817 -0.080 5.079 0.080 ;
      RECT 4.727 -0.080 4.817 0.122 ;
      RECT 4.037 -0.080 4.727 0.080 ;
      RECT 3.947 -0.080 4.037 0.370 ;
      RECT 3.422 -0.080 3.947 0.080 ;
      RECT 3.332 -0.080 3.422 0.287 ;
      RECT 2.741 -0.080 3.332 0.080 ;
      RECT 2.651 -0.080 2.741 0.122 ;
      RECT 1.828 -0.080 2.651 0.080 ;
      RECT 1.738 -0.080 1.828 0.122 ;
      RECT 1.118 -0.080 1.738 0.080 ;
      RECT 1.028 -0.080 1.118 0.122 ;
      RECT 0.296 -0.080 1.028 0.080 ;
      RECT 0.206 -0.080 0.296 0.122 ;
      RECT 0.000 -0.080 0.206 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.194 1.120 5.400 1.280 ;
      RECT 5.081 1.078 5.194 1.280 ;
      RECT 4.806 1.120 5.081 1.280 ;
      RECT 4.716 1.078 4.806 1.280 ;
      RECT 3.250 1.120 4.716 1.280 ;
      RECT 3.161 1.078 3.250 1.280 ;
      RECT 2.695 1.120 3.161 1.280 ;
      RECT 2.634 0.902 2.695 1.280 ;
      RECT 1.824 1.120 2.634 1.280 ;
      RECT 1.734 1.078 1.824 1.280 ;
      RECT 1.115 1.120 1.734 1.280 ;
      RECT 1.025 1.078 1.115 1.280 ;
      RECT 0.311 1.120 1.025 1.280 ;
      RECT 0.222 1.078 0.311 1.280 ;
      RECT 0.000 1.120 0.222 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.124 0.500 5.214 0.581 ;
      RECT 4.994 0.513 5.124 0.568 ;
      RECT 4.994 0.742 5.008 0.935 ;
      RECT 4.984 0.513 4.994 0.935 ;
      RECT 4.924 0.307 4.984 0.935 ;
      RECT 4.895 0.307 4.924 0.388 ;
      RECT 4.918 0.742 4.924 0.935 ;
      RECT 4.707 0.855 4.918 0.910 ;
      RECT 4.757 0.524 4.847 0.605 ;
      RECT 4.679 0.524 4.757 0.579 ;
      RECT 4.707 0.683 4.722 0.764 ;
      RECT 4.646 0.683 4.707 0.910 ;
      RECT 4.664 0.480 4.679 0.579 ;
      RECT 4.603 0.151 4.664 0.579 ;
      RECT 4.632 0.683 4.646 0.764 ;
      RECT 4.455 0.855 4.646 0.910 ;
      RECT 4.402 0.151 4.603 0.206 ;
      RECT 4.464 0.480 4.603 0.535 ;
      RECT 4.482 0.298 4.542 0.387 ;
      RECT 4.339 0.332 4.482 0.387 ;
      RECT 4.455 0.480 4.464 0.771 ;
      RECT 4.404 0.480 4.455 0.800 ;
      RECT 4.394 0.855 4.455 1.050 ;
      RECT 4.394 0.717 4.404 0.800 ;
      RECT 4.342 0.151 4.402 0.268 ;
      RECT 3.373 0.995 4.394 1.050 ;
      RECT 4.334 0.332 4.339 0.669 ;
      RECT 4.278 0.332 4.334 0.940 ;
      RECT 4.273 0.614 4.278 0.940 ;
      RECT 3.496 0.886 4.273 0.940 ;
      RECT 4.152 0.271 4.212 0.780 ;
      RECT 4.025 0.508 4.086 0.831 ;
      RECT 3.618 0.776 4.025 0.831 ;
      RECT 3.760 0.665 3.847 0.720 ;
      RECT 3.760 0.317 3.826 0.371 ;
      RECT 3.699 0.150 3.760 0.720 ;
      RECT 3.558 0.233 3.618 0.831 ;
      RECT 3.245 0.554 3.558 0.608 ;
      RECT 3.435 0.843 3.496 0.940 ;
      RECT 3.431 0.357 3.492 0.462 ;
      RECT 2.938 0.843 3.435 0.898 ;
      RECT 3.102 0.357 3.431 0.412 ;
      RECT 3.312 0.954 3.373 1.050 ;
      RECT 2.816 0.954 3.312 1.008 ;
      RECT 3.059 0.244 3.102 0.650 ;
      RECT 3.042 0.244 3.059 0.783 ;
      RECT 2.973 0.244 3.042 0.299 ;
      RECT 2.998 0.595 3.042 0.783 ;
      RECT 2.759 0.394 2.965 0.449 ;
      RECT 2.877 0.665 2.938 0.898 ;
      RECT 2.759 0.665 2.877 0.720 ;
      RECT 2.755 0.776 2.816 1.008 ;
      RECT 2.699 0.257 2.759 0.720 ;
      RECT 2.336 0.776 2.755 0.831 ;
      RECT 2.535 0.257 2.699 0.312 ;
      RECT 2.419 0.665 2.699 0.720 ;
      RECT 2.445 0.231 2.535 0.312 ;
      RECT 1.979 0.982 2.449 1.037 ;
      RECT 2.275 0.306 2.336 0.915 ;
      RECT 2.146 0.390 2.199 0.902 ;
      RECT 2.138 0.306 2.146 0.902 ;
      RECT 2.085 0.306 2.138 0.445 ;
      RECT 2.071 0.833 2.138 0.902 ;
      RECT 2.024 0.542 2.076 0.631 ;
      RECT 1.441 0.833 2.071 0.888 ;
      RECT 2.024 0.150 2.060 0.205 ;
      RECT 1.964 0.150 2.024 0.749 ;
      RECT 1.919 0.954 1.979 1.037 ;
      RECT 1.618 0.192 1.964 0.246 ;
      RECT 0.672 0.954 1.919 1.008 ;
      RECT 1.837 0.375 1.898 0.482 ;
      RECT 1.618 0.427 1.837 0.482 ;
      RECT 1.618 0.681 1.661 0.736 ;
      RECT 1.618 0.302 1.654 0.357 ;
      RECT 1.557 0.161 1.618 0.246 ;
      RECT 1.557 0.302 1.618 0.736 ;
      RECT 1.302 0.161 1.557 0.215 ;
      RECT 1.526 0.526 1.557 0.613 ;
      RECT 1.380 0.287 1.441 0.888 ;
      RECT 1.011 0.833 1.380 0.888 ;
      RECT 1.246 0.300 1.306 0.725 ;
      RECT 1.176 0.300 1.246 0.355 ;
      RECT 1.176 0.670 1.246 0.725 ;
      RECT 0.950 0.202 1.011 0.888 ;
      RECT 0.892 0.202 0.950 0.257 ;
      RECT 0.800 0.833 0.950 0.888 ;
      RECT 0.831 0.163 0.892 0.257 ;
      RECT 0.827 0.318 0.888 0.733 ;
      RECT 0.800 0.163 0.831 0.218 ;
      RECT 0.788 0.469 0.827 0.554 ;
      RECT 0.672 0.343 0.703 0.501 ;
      RECT 0.643 0.343 0.672 1.008 ;
      RECT 0.611 0.446 0.643 1.008 ;
      RECT 0.471 0.935 0.532 1.050 ;
      RECT 0.478 0.343 0.507 0.424 ;
      RECT 0.478 0.746 0.486 0.827 ;
      RECT 0.417 0.343 0.478 0.827 ;
      RECT 0.137 0.935 0.471 0.989 ;
      RECT 0.396 0.746 0.417 0.827 ;
      RECT 0.108 0.343 0.137 0.424 ;
      RECT 0.108 0.746 0.137 0.989 ;
      RECT 0.077 0.343 0.108 0.989 ;
      RECT 0.048 0.343 0.077 0.827 ;
  END
END SEDFFHQX1

MACRO SDFFSHQXL
  CLASS CORE ;
  FOREIGN SDFFSHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.618 0.521 3.698 0.602 ;
      RECT 3.607 0.521 3.618 0.627 ;
      RECT 3.578 0.529 3.607 0.627 ;
      RECT 3.517 0.529 3.578 0.994 ;
      RECT 2.136 0.939 3.517 0.994 ;
      RECT 2.075 0.633 2.136 0.994 ;
      RECT 2.043 0.633 2.075 0.701 ;
      RECT 1.982 0.573 2.043 0.701 ;
      RECT 1.804 0.608 1.982 0.701 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.757 0.435 0.864 0.535 ;
      RECT 0.688 0.480 0.757 0.535 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.882 0.590 0.943 0.781 ;
      RECT 0.818 0.700 0.882 0.781 ;
      RECT 0.643 0.726 0.818 0.781 ;
      RECT 0.616 0.706 0.643 0.781 ;
      RECT 0.555 0.614 0.616 0.781 ;
      RECT 0.408 0.614 0.555 0.669 ;
      RECT 0.347 0.579 0.408 0.669 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.082 0.267 4.143 0.715 ;
      RECT 4.013 0.267 4.082 0.348 ;
      RECT 4.062 0.627 4.082 0.715 ;
      RECT 3.835 0.661 4.062 0.715 ;
      RECT 3.774 0.661 3.835 0.824 ;
      RECT 3.745 0.743 3.774 0.824 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.168 0.351 1.172 0.465 ;
      RECT 1.107 0.351 1.168 0.494 ;
      RECT 1.054 0.351 1.107 0.485 ;
      RECT 1.031 0.351 1.054 0.465 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.137 0.211 0.139 0.292 ;
      RECT 0.034 0.162 0.137 0.292 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.764 -0.080 4.200 0.080 ;
      RECT 3.674 -0.080 3.764 0.325 ;
      RECT 3.312 -0.080 3.674 0.080 ;
      RECT 3.222 -0.080 3.312 0.122 ;
      RECT 2.520 -0.080 3.222 0.080 ;
      RECT 2.459 -0.080 2.520 0.341 ;
      RECT 1.771 -0.080 2.459 0.080 ;
      RECT 1.681 -0.080 1.771 0.186 ;
      RECT 0.843 -0.080 1.681 0.080 ;
      RECT 0.753 -0.080 0.843 0.122 ;
      RECT 0.297 -0.080 0.753 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.026 1.120 4.200 1.280 ;
      RECT 3.936 0.805 4.026 1.280 ;
      RECT 3.674 1.120 3.936 1.280 ;
      RECT 3.584 1.078 3.674 1.280 ;
      RECT 3.308 1.120 3.584 1.280 ;
      RECT 3.218 1.078 3.308 1.280 ;
      RECT 2.466 1.120 3.218 1.280 ;
      RECT 2.369 1.078 2.466 1.280 ;
      RECT 2.013 1.120 2.369 1.280 ;
      RECT 1.763 1.001 2.013 1.280 ;
      RECT 0.902 1.120 1.763 1.280 ;
      RECT 0.811 1.078 0.902 1.280 ;
      RECT 0.292 1.120 0.811 1.280 ;
      RECT 0.202 1.078 0.292 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.998 0.515 4.000 0.583 ;
      RECT 3.939 0.411 3.998 0.583 ;
      RECT 3.938 0.411 3.939 0.570 ;
      RECT 3.512 0.411 3.938 0.465 ;
      RECT 3.481 0.192 3.512 0.465 ;
      RECT 3.451 0.165 3.481 0.465 ;
      RECT 3.387 0.165 3.451 0.248 ;
      RECT 3.389 0.629 3.443 0.750 ;
      RECT 3.382 0.307 3.389 0.750 ;
      RECT 3.235 0.193 3.387 0.248 ;
      RECT 3.328 0.307 3.382 0.683 ;
      RECT 3.153 0.629 3.328 0.683 ;
      RECT 3.174 0.193 3.235 0.539 ;
      RECT 2.950 0.193 3.174 0.248 ;
      RECT 3.031 0.485 3.174 0.539 ;
      RECT 3.092 0.629 3.153 0.714 ;
      RECT 2.970 0.340 3.060 0.421 ;
      RECT 2.483 0.819 3.051 0.874 ;
      RECT 2.970 0.485 3.031 0.760 ;
      RECT 2.909 0.367 2.970 0.421 ;
      RECT 2.800 0.705 2.970 0.760 ;
      RECT 2.860 0.180 2.950 0.261 ;
      RECT 2.848 0.367 2.909 0.582 ;
      RECT 2.744 0.527 2.848 0.582 ;
      RECT 2.719 0.263 2.748 0.344 ;
      RECT 2.683 0.527 2.744 0.614 ;
      RECT 2.658 0.263 2.719 0.468 ;
      RECT 2.618 0.705 2.665 0.760 ;
      RECT 2.618 0.413 2.658 0.468 ;
      RECT 2.557 0.413 2.618 0.760 ;
      RECT 2.422 0.445 2.483 0.874 ;
      RECT 2.396 0.445 2.422 0.500 ;
      RECT 2.390 0.808 2.422 0.874 ;
      RECT 2.335 0.321 2.396 0.500 ;
      RECT 2.287 0.808 2.390 0.863 ;
      RECT 2.274 0.555 2.360 0.636 ;
      RECT 2.308 0.321 2.335 0.376 ;
      RECT 2.247 0.161 2.308 0.376 ;
      RECT 2.197 0.795 2.287 0.876 ;
      RECT 2.270 0.431 2.274 0.636 ;
      RECT 2.213 0.431 2.270 0.623 ;
      RECT 2.158 0.161 2.247 0.215 ;
      RECT 2.172 0.431 2.213 0.486 ;
      RECT 2.111 0.318 2.172 0.486 ;
      RECT 2.015 0.318 2.111 0.475 ;
      RECT 1.926 0.185 2.043 0.239 ;
      RECT 1.743 0.420 2.015 0.475 ;
      RECT 1.743 0.808 1.936 0.863 ;
      RECT 1.865 0.185 1.926 0.325 ;
      RECT 1.493 0.270 1.865 0.325 ;
      RECT 1.682 0.420 1.743 0.863 ;
      RECT 1.579 0.449 1.682 0.504 ;
      RECT 1.560 0.562 1.621 0.865 ;
      RECT 1.491 0.562 1.560 0.617 ;
      RECT 1.436 0.811 1.560 0.865 ;
      RECT 1.320 0.673 1.499 0.727 ;
      RECT 1.491 0.242 1.493 0.325 ;
      RECT 1.430 0.242 1.491 0.617 ;
      RECT 1.346 0.811 1.436 0.892 ;
      RECT 1.319 0.242 1.430 0.296 ;
      RECT 1.259 0.365 1.320 0.727 ;
      RECT 1.092 0.673 1.259 0.727 ;
      RECT 1.156 0.845 1.217 1.007 ;
      RECT 1.104 0.171 1.195 0.252 ;
      RECT 0.438 0.952 1.156 1.007 ;
      RECT 0.468 0.194 1.104 0.249 ;
      RECT 1.031 0.673 1.092 0.896 ;
      RECT 0.138 0.842 1.031 0.896 ;
      RECT 0.537 0.318 0.939 0.373 ;
      RECT 0.537 0.452 0.586 0.557 ;
      RECT 0.525 0.318 0.537 0.557 ;
      RECT 0.476 0.318 0.525 0.524 ;
      RECT 0.261 0.732 0.495 0.787 ;
      RECT 0.445 0.346 0.476 0.524 ;
      RECT 0.407 0.152 0.468 0.249 ;
      RECT 0.261 0.469 0.445 0.524 ;
      RECT 0.200 0.469 0.261 0.787 ;
      RECT 0.098 0.750 0.138 0.896 ;
      RECT 0.098 0.346 0.123 0.456 ;
      RECT 0.077 0.346 0.098 0.896 ;
      RECT 0.062 0.346 0.077 0.831 ;
      RECT 0.048 0.401 0.062 0.831 ;
      RECT 0.037 0.401 0.048 0.807 ;
  END
END SDFFSHQXL

MACRO SDFFSHQX4
  CLASS CORE ;
  FOREIGN SDFFSHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.132 0.536 5.192 0.590 ;
      RECT 5.043 0.536 5.132 0.611 ;
      RECT 4.692 0.556 5.043 0.611 ;
      RECT 4.680 0.537 4.692 0.611 ;
      RECT 4.619 0.537 4.680 1.008 ;
      RECT 4.582 0.537 4.619 0.592 ;
      RECT 4.587 0.894 4.619 1.008 ;
      RECT 3.363 0.954 4.587 1.008 ;
      RECT 3.302 0.840 3.363 1.008 ;
      RECT 2.197 0.840 3.302 0.895 ;
      RECT 2.197 0.706 2.218 0.761 ;
      RECT 2.136 0.690 2.197 0.895 ;
      RECT 1.875 0.690 2.136 0.745 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.818 0.595 0.837 0.676 ;
      RECT 0.757 0.321 0.818 0.676 ;
      RECT 0.721 0.321 0.757 0.376 ;
      RECT 0.746 0.595 0.757 0.676 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.456 0.573 0.468 0.646 ;
      RECT 0.334 0.567 0.456 0.669 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.547 0.190 5.552 0.306 ;
      RECT 5.486 0.190 5.547 0.758 ;
      RECT 5.462 0.190 5.486 0.356 ;
      RECT 5.388 0.704 5.486 0.758 ;
      RECT 4.873 0.301 5.462 0.356 ;
      RECT 5.287 0.700 5.388 1.033 ;
      RECT 5.229 0.711 5.287 0.960 ;
      RECT 5.193 0.711 5.229 0.767 ;
      RECT 4.957 0.711 5.193 0.765 ;
      RECT 4.916 0.711 4.957 0.767 ;
      RECT 4.826 0.711 4.916 0.935 ;
      RECT 4.811 0.251 4.873 0.356 ;
      RECT 4.783 0.251 4.811 0.332 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.077 0.329 1.188 0.500 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.245 0.418 0.331 0.510 ;
      RECT 0.184 0.418 0.245 0.555 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.213 -0.080 5.600 0.080 ;
      RECT 5.123 -0.080 5.213 0.212 ;
      RECT 4.173 -0.080 5.123 0.080 ;
      RECT 4.083 -0.080 4.173 0.122 ;
      RECT 3.039 -0.080 4.083 0.080 ;
      RECT 2.948 -0.080 3.039 0.290 ;
      RECT 2.655 -0.080 2.948 0.080 ;
      RECT 2.565 -0.080 2.655 0.317 ;
      RECT 1.783 -0.080 2.565 0.080 ;
      RECT 1.693 -0.080 1.783 0.233 ;
      RECT 0.912 -0.080 1.693 0.080 ;
      RECT 0.822 -0.080 0.912 0.122 ;
      RECT 0.343 -0.080 0.822 0.080 ;
      RECT 0.253 -0.080 0.343 0.122 ;
      RECT 0.000 -0.080 0.253 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.530 1.120 5.600 1.280 ;
      RECT 5.469 0.844 5.530 1.280 ;
      RECT 5.117 1.120 5.469 1.280 ;
      RECT 5.027 0.844 5.117 1.280 ;
      RECT 4.704 1.120 5.027 1.280 ;
      RECT 4.614 1.078 4.704 1.280 ;
      RECT 4.314 1.120 4.614 1.280 ;
      RECT 4.224 1.078 4.314 1.280 ;
      RECT 3.073 1.120 4.224 1.280 ;
      RECT 2.983 1.078 3.073 1.280 ;
      RECT 2.669 1.120 2.983 1.280 ;
      RECT 2.579 1.078 2.669 1.280 ;
      RECT 2.280 1.120 2.579 1.280 ;
      RECT 2.190 1.078 2.280 1.280 ;
      RECT 1.877 1.120 2.190 1.280 ;
      RECT 1.787 1.078 1.877 1.280 ;
      RECT 1.009 1.120 1.787 1.280 ;
      RECT 0.919 1.004 1.009 1.280 ;
      RECT 0.345 1.120 0.919 1.280 ;
      RECT 0.255 1.078 0.345 1.280 ;
      RECT 0.000 1.120 0.255 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.396 0.525 5.425 0.606 ;
      RECT 5.335 0.424 5.396 0.606 ;
      RECT 4.964 0.424 5.335 0.479 ;
      RECT 4.858 0.424 4.964 0.492 ;
      RECT 4.681 0.424 4.858 0.479 ;
      RECT 4.620 0.206 4.681 0.479 ;
      RECT 3.936 0.206 4.620 0.261 ;
      RECT 4.494 0.714 4.523 0.795 ;
      RECT 4.433 0.368 4.494 0.795 ;
      RECT 4.216 0.368 4.433 0.423 ;
      RECT 4.334 0.536 4.363 0.617 ;
      RECT 4.273 0.536 4.334 0.899 ;
      RECT 3.936 0.844 4.273 0.899 ;
      RECT 4.126 0.336 4.216 0.423 ;
      RECT 4.116 0.367 4.126 0.423 ;
      RECT 4.041 0.367 4.116 0.558 ;
      RECT 4.026 0.477 4.041 0.558 ;
      RECT 3.875 0.206 3.936 0.899 ;
      RECT 3.802 0.206 3.875 0.261 ;
      RECT 3.463 0.844 3.875 0.899 ;
      RECT 3.773 0.206 3.802 0.336 ;
      RECT 3.712 0.173 3.773 0.336 ;
      RECT 3.585 0.731 3.755 0.786 ;
      RECT 3.420 0.173 3.712 0.227 ;
      RECT 3.585 0.286 3.611 0.367 ;
      RECT 3.524 0.286 3.585 0.786 ;
      RECT 3.521 0.286 3.524 0.415 ;
      RECT 3.253 0.731 3.524 0.786 ;
      RECT 3.230 0.361 3.521 0.415 ;
      RECT 3.359 0.173 3.420 0.304 ;
      RECT 3.330 0.223 3.359 0.304 ;
      RECT 2.637 0.470 3.358 0.525 ;
      RECT 3.192 0.711 3.253 0.786 ;
      RECT 3.139 0.262 3.230 0.415 ;
      RECT 3.154 0.951 3.215 1.049 ;
      RECT 2.870 0.711 3.192 0.765 ;
      RECT 1.627 0.951 3.154 1.006 ;
      RECT 2.848 0.361 3.139 0.415 ;
      RECT 2.780 0.685 2.870 0.765 ;
      RECT 2.772 0.264 2.848 0.415 ;
      RECT 2.758 0.264 2.772 0.345 ;
      RECT 2.576 0.430 2.637 0.751 ;
      RECT 2.446 0.430 2.576 0.485 ;
      RECT 2.504 0.683 2.576 0.751 ;
      RECT 2.194 0.546 2.511 0.601 ;
      RECT 2.414 0.683 2.504 0.764 ;
      RECT 2.385 0.185 2.446 0.485 ;
      RECT 1.986 0.185 2.385 0.239 ;
      RECT 2.176 0.310 2.194 0.635 ;
      RECT 2.133 0.296 2.176 0.635 ;
      RECT 2.085 0.296 2.133 0.377 ;
      RECT 1.725 0.580 2.133 0.635 ;
      RECT 1.548 0.470 2.072 0.525 ;
      RECT 2.003 0.801 2.064 0.895 ;
      RECT 1.725 0.801 2.003 0.856 ;
      RECT 1.925 0.185 1.986 0.406 ;
      RECT 1.624 0.351 1.925 0.406 ;
      RECT 1.664 0.580 1.725 0.856 ;
      RECT 1.551 0.951 1.627 1.008 ;
      RECT 1.563 0.151 1.624 0.406 ;
      RECT 1.515 0.151 1.563 0.206 ;
      RECT 1.425 0.954 1.551 1.008 ;
      RECT 1.487 0.470 1.548 0.885 ;
      RECT 1.454 0.470 1.487 0.525 ;
      RECT 1.393 0.198 1.454 0.525 ;
      RECT 1.364 0.732 1.425 1.008 ;
      RECT 1.363 0.198 1.393 0.252 ;
      RECT 1.330 0.732 1.364 0.787 ;
      RECT 1.269 0.346 1.330 0.787 ;
      RECT 1.226 0.856 1.287 0.964 ;
      RECT 0.733 0.732 1.269 0.787 ;
      RECT 0.541 0.194 1.262 0.249 ;
      RECT 0.856 0.856 1.226 0.911 ;
      RECT 0.795 0.856 0.856 1.023 ;
      RECT 0.514 0.968 0.795 1.023 ;
      RECT 0.672 0.732 0.733 0.913 ;
      RECT 0.141 0.858 0.672 0.913 ;
      RECT 0.610 0.493 0.640 0.574 ;
      RECT 0.549 0.374 0.610 0.789 ;
      RECT 0.545 0.374 0.549 0.429 ;
      RECT 0.430 0.735 0.549 0.789 ;
      RECT 0.455 0.348 0.545 0.429 ;
      RECT 0.465 0.155 0.541 0.249 ;
      RECT 0.451 0.155 0.465 0.236 ;
      RECT 0.111 0.281 0.141 0.362 ;
      RECT 0.111 0.714 0.141 0.938 ;
      RECT 0.050 0.281 0.111 0.938 ;
  END
END SDFFSHQX4

MACRO SDFFSHQX2
  CLASS CORE ;
  FOREIGN SDFFSHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.652 0.502 4.713 0.894 ;
      RECT 4.071 0.839 4.652 0.894 ;
      RECT 4.071 0.518 4.089 0.599 ;
      RECT 4.010 0.518 4.071 0.894 ;
      RECT 3.998 0.518 4.010 0.599 ;
      RECT 3.991 0.839 4.010 0.894 ;
      RECT 3.930 0.839 3.991 1.025 ;
      RECT 2.917 0.970 3.930 1.025 ;
      RECT 2.856 0.870 2.917 1.025 ;
      RECT 2.837 0.870 2.856 0.973 ;
      RECT 2.588 0.870 2.837 0.925 ;
      RECT 2.537 0.870 2.588 0.973 ;
      RECT 2.477 0.870 2.537 1.039 ;
      RECT 2.064 0.985 2.477 1.039 ;
      RECT 2.043 0.585 2.064 1.039 ;
      RECT 2.003 0.573 2.043 1.039 ;
      RECT 1.791 0.573 2.003 0.639 ;
      RECT 1.716 0.573 1.791 0.662 ;
      RECT 1.701 0.581 1.716 0.662 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.693 0.548 0.831 0.657 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.346 0.485 0.427 0.565 ;
      RECT 0.337 0.444 0.346 0.565 ;
      RECT 0.293 0.444 0.337 0.552 ;
      RECT 0.285 0.439 0.293 0.552 ;
      RECT 0.232 0.439 0.285 0.499 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.522 0.307 4.583 0.733 ;
      RECT 4.493 0.307 4.522 0.367 ;
      RECT 4.432 0.679 4.522 0.733 ;
      RECT 4.468 0.307 4.493 0.362 ;
      RECT 4.378 0.281 4.468 0.362 ;
      RECT 4.343 0.679 4.432 0.760 ;
      RECT 4.257 0.679 4.343 0.761 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.945 0.435 1.057 0.557 ;
      RECT 0.932 0.439 0.945 0.494 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.126 0.906 0.179 1.008 ;
      RECT 0.057 0.906 0.126 1.027 ;
      RECT 0.050 0.906 0.057 1.008 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.807 -0.080 4.900 0.080 ;
      RECT 4.717 -0.080 4.807 0.345 ;
      RECT 3.830 -0.080 4.717 0.080 ;
      RECT 3.740 -0.080 3.830 0.122 ;
      RECT 2.897 -0.080 3.740 0.080 ;
      RECT 2.807 -0.080 2.897 0.303 ;
      RECT 2.500 -0.080 2.807 0.080 ;
      RECT 2.439 -0.080 2.500 0.311 ;
      RECT 1.725 -0.080 2.439 0.080 ;
      RECT 1.635 -0.080 1.725 0.214 ;
      RECT 0.833 -0.080 1.635 0.080 ;
      RECT 0.742 -0.080 0.833 0.122 ;
      RECT 0.286 -0.080 0.742 0.080 ;
      RECT 0.196 -0.080 0.286 0.122 ;
      RECT 0.000 -0.080 0.196 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.549 1.120 4.900 1.280 ;
      RECT 4.459 0.988 4.549 1.280 ;
      RECT 4.151 1.120 4.459 1.280 ;
      RECT 4.061 0.976 4.151 1.280 ;
      RECT 2.755 1.120 4.061 1.280 ;
      RECT 2.665 0.996 2.755 1.280 ;
      RECT 1.942 1.120 2.665 1.280 ;
      RECT 1.727 1.001 1.942 1.280 ;
      RECT 0.895 1.120 1.727 1.280 ;
      RECT 0.805 1.001 0.895 1.280 ;
      RECT 0.289 1.120 0.805 1.280 ;
      RECT 0.199 1.078 0.289 1.280 ;
      RECT 0.000 1.120 0.199 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.213 0.499 4.429 0.554 ;
      RECT 4.152 0.206 4.213 0.554 ;
      RECT 3.477 0.206 4.152 0.261 ;
      RECT 3.821 0.506 3.869 0.892 ;
      RECT 3.808 0.506 3.821 0.905 ;
      RECT 3.788 0.506 3.808 0.561 ;
      RECT 3.731 0.824 3.808 0.905 ;
      RECT 3.788 0.348 3.802 0.429 ;
      RECT 3.727 0.348 3.788 0.561 ;
      RECT 3.655 0.657 3.745 0.738 ;
      RECT 3.712 0.348 3.727 0.429 ;
      RECT 3.723 0.490 3.727 0.561 ;
      RECT 3.633 0.490 3.723 0.571 ;
      RECT 3.477 0.670 3.655 0.725 ;
      RECT 3.435 0.206 3.477 0.915 ;
      RECT 3.416 0.189 3.435 0.915 ;
      RECT 3.374 0.189 3.416 0.381 ;
      RECT 3.057 0.861 3.416 0.915 ;
      RECT 3.082 0.189 3.374 0.244 ;
      RECT 3.287 0.746 3.354 0.801 ;
      RECT 3.273 0.380 3.287 0.801 ;
      RECT 3.226 0.305 3.273 0.801 ;
      RECT 3.183 0.305 3.226 0.435 ;
      RECT 2.956 0.746 3.226 0.801 ;
      RECT 2.706 0.380 3.183 0.435 ;
      RECT 2.414 0.489 3.162 0.544 ;
      RECT 3.021 0.189 3.082 0.325 ;
      RECT 2.992 0.244 3.021 0.325 ;
      RECT 2.866 0.733 2.956 0.814 ;
      RECT 2.565 0.746 2.866 0.801 ;
      RECT 2.645 0.265 2.706 0.435 ;
      RECT 2.616 0.265 2.645 0.346 ;
      RECT 2.475 0.733 2.565 0.814 ;
      RECT 2.353 0.417 2.414 0.915 ;
      RECT 2.315 0.417 2.353 0.471 ;
      RECT 2.305 0.835 2.353 0.915 ;
      RECT 2.288 0.336 2.315 0.471 ;
      RECT 2.250 0.848 2.305 0.915 ;
      RECT 2.254 0.161 2.288 0.471 ;
      RECT 2.225 0.533 2.286 0.685 ;
      RECT 2.227 0.161 2.254 0.390 ;
      RECT 2.160 0.848 2.250 0.929 ;
      RECT 2.117 0.161 2.227 0.215 ;
      RECT 2.190 0.533 2.225 0.588 ;
      RECT 2.129 0.446 2.190 0.588 ;
      RECT 2.091 0.446 2.129 0.501 ;
      RECT 2.030 0.337 2.091 0.501 ;
      RECT 2.001 0.337 2.030 0.449 ;
      RECT 1.937 0.171 2.027 0.252 ;
      RECT 1.598 0.394 2.001 0.449 ;
      RECT 1.905 0.198 1.937 0.252 ;
      RECT 1.844 0.198 1.905 0.338 ;
      RECT 1.808 0.779 1.898 0.860 ;
      RECT 1.384 0.283 1.844 0.338 ;
      RECT 1.598 0.792 1.808 0.846 ;
      RECT 1.598 0.517 1.612 0.598 ;
      RECT 1.537 0.394 1.598 0.846 ;
      RECT 1.522 0.517 1.537 0.598 ;
      RECT 1.399 0.930 1.489 1.011 ;
      RECT 1.262 0.943 1.399 0.998 ;
      RECT 1.323 0.283 1.384 0.850 ;
      RECT 1.267 0.323 1.323 0.377 ;
      RECT 1.233 0.732 1.262 0.998 ;
      RECT 1.233 0.442 1.248 0.523 ;
      RECT 1.201 0.442 1.233 0.998 ;
      RECT 1.173 0.156 1.209 0.211 ;
      RECT 1.172 0.442 1.201 0.787 ;
      RECT 1.112 0.156 1.173 0.261 ;
      RECT 1.157 0.442 1.172 0.523 ;
      RECT 0.595 0.732 1.172 0.787 ;
      RECT 1.079 0.856 1.140 0.979 ;
      RECT 0.472 0.206 1.112 0.261 ;
      RECT 0.729 0.856 1.079 0.911 ;
      RECT 0.593 0.315 0.920 0.370 ;
      RECT 0.668 0.856 0.729 1.023 ;
      RECT 0.443 0.968 0.668 1.023 ;
      RECT 0.534 0.732 0.595 0.913 ;
      RECT 0.532 0.315 0.593 0.677 ;
      RECT 0.350 0.858 0.534 0.913 ;
      RECT 0.526 0.315 0.532 0.424 ;
      RECT 0.473 0.623 0.532 0.677 ;
      RECT 0.408 0.343 0.526 0.424 ;
      RECT 0.412 0.623 0.473 0.779 ;
      RECT 0.411 0.150 0.472 0.261 ;
      RECT 0.382 0.150 0.411 0.231 ;
      RECT 0.289 0.773 0.350 0.913 ;
      RECT 0.138 0.773 0.289 0.827 ;
      RECT 0.099 0.323 0.138 0.404 ;
      RECT 0.099 0.746 0.138 0.827 ;
      RECT 0.048 0.323 0.099 0.827 ;
      RECT 0.038 0.349 0.048 0.814 ;
  END
END SDFFSHQX2

MACRO SDFFSHQX1
  CLASS CORE ;
  FOREIGN SDFFSHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.732 0.439 3.793 0.500 ;
      RECT 3.698 0.445 3.732 0.500 ;
      RECT 3.637 0.445 3.698 0.583 ;
      RECT 3.607 0.502 3.637 0.583 ;
      RECT 3.578 0.529 3.607 0.583 ;
      RECT 3.517 0.529 3.578 0.994 ;
      RECT 2.136 0.939 3.517 0.994 ;
      RECT 2.075 0.633 2.136 0.994 ;
      RECT 2.043 0.633 2.075 0.701 ;
      RECT 1.982 0.573 2.043 0.701 ;
      RECT 1.804 0.608 1.982 0.701 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.810 0.344 0.818 0.661 ;
      RECT 0.793 0.344 0.810 0.674 ;
      RECT 0.757 0.331 0.793 0.674 ;
      RECT 0.737 0.331 0.757 0.439 ;
      RECT 0.720 0.593 0.757 0.674 ;
      RECT 0.703 0.331 0.737 0.412 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.374 0.539 0.496 0.669 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.082 0.204 4.143 0.715 ;
      RECT 4.062 0.204 4.082 0.307 ;
      RECT 4.062 0.627 4.082 0.715 ;
      RECT 4.028 0.204 4.062 0.290 ;
      RECT 3.835 0.661 4.062 0.715 ;
      RECT 3.774 0.661 3.835 0.819 ;
      RECT 3.745 0.738 3.774 0.819 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.031 0.421 1.172 0.536 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.273 0.439 0.293 0.494 ;
      RECT 0.269 0.439 0.273 0.565 ;
      RECT 0.221 0.439 0.269 0.567 ;
      RECT 0.208 0.439 0.221 0.598 ;
      RECT 0.160 0.511 0.208 0.598 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.753 -0.080 4.200 0.080 ;
      RECT 3.663 -0.080 3.753 0.122 ;
      RECT 3.312 -0.080 3.663 0.080 ;
      RECT 3.222 -0.080 3.312 0.122 ;
      RECT 2.520 -0.080 3.222 0.080 ;
      RECT 2.459 -0.080 2.520 0.290 ;
      RECT 1.771 -0.080 2.459 0.080 ;
      RECT 1.681 -0.080 1.771 0.186 ;
      RECT 0.835 -0.080 1.681 0.080 ;
      RECT 0.745 -0.080 0.835 0.122 ;
      RECT 0.286 -0.080 0.745 0.080 ;
      RECT 0.196 -0.080 0.286 0.206 ;
      RECT 0.000 -0.080 0.196 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.026 1.120 4.200 1.280 ;
      RECT 3.936 0.805 4.026 1.280 ;
      RECT 3.680 1.120 3.936 1.280 ;
      RECT 3.590 1.078 3.680 1.280 ;
      RECT 3.308 1.120 3.590 1.280 ;
      RECT 3.218 1.078 3.308 1.280 ;
      RECT 2.466 1.120 3.218 1.280 ;
      RECT 2.369 1.078 2.466 1.280 ;
      RECT 2.013 1.120 2.369 1.280 ;
      RECT 1.763 1.001 2.013 1.280 ;
      RECT 0.986 1.120 1.763 1.280 ;
      RECT 0.925 1.002 0.986 1.280 ;
      RECT 0.292 1.120 0.925 1.280 ;
      RECT 0.202 1.078 0.292 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.964 0.502 3.993 0.583 ;
      RECT 3.903 0.306 3.964 0.583 ;
      RECT 3.512 0.306 3.903 0.361 ;
      RECT 3.481 0.192 3.512 0.361 ;
      RECT 3.451 0.165 3.481 0.361 ;
      RECT 3.393 0.629 3.454 0.750 ;
      RECT 3.387 0.165 3.451 0.246 ;
      RECT 3.389 0.629 3.393 0.683 ;
      RECT 3.328 0.314 3.389 0.683 ;
      RECT 3.187 0.192 3.387 0.246 ;
      RECT 3.167 0.629 3.328 0.683 ;
      RECT 3.126 0.192 3.187 0.539 ;
      RECT 3.077 0.629 3.167 0.710 ;
      RECT 2.998 0.192 3.126 0.246 ;
      RECT 2.972 0.485 3.126 0.539 ;
      RECT 2.848 0.345 3.060 0.400 ;
      RECT 2.483 0.819 3.051 0.874 ;
      RECT 2.935 0.192 2.998 0.290 ;
      RECT 2.911 0.485 2.972 0.760 ;
      RECT 2.828 0.236 2.935 0.290 ;
      RECT 2.800 0.705 2.911 0.760 ;
      RECT 2.787 0.345 2.848 0.582 ;
      RECT 2.744 0.527 2.787 0.582 ;
      RECT 2.683 0.527 2.744 0.614 ;
      RECT 2.697 0.257 2.726 0.338 ;
      RECT 2.636 0.257 2.697 0.437 ;
      RECT 2.618 0.705 2.677 0.760 ;
      RECT 2.618 0.382 2.636 0.437 ;
      RECT 2.557 0.382 2.618 0.760 ;
      RECT 2.422 0.380 2.483 0.874 ;
      RECT 2.396 0.380 2.422 0.435 ;
      RECT 2.390 0.804 2.422 0.874 ;
      RECT 2.335 0.321 2.396 0.435 ;
      RECT 2.287 0.804 2.390 0.871 ;
      RECT 2.274 0.561 2.360 0.615 ;
      RECT 2.323 0.321 2.335 0.376 ;
      RECT 2.294 0.295 2.323 0.376 ;
      RECT 2.248 0.163 2.294 0.376 ;
      RECT 2.197 0.790 2.287 0.871 ;
      RECT 2.213 0.431 2.274 0.615 ;
      RECT 2.233 0.150 2.248 0.376 ;
      RECT 2.158 0.150 2.233 0.231 ;
      RECT 2.141 0.431 2.213 0.486 ;
      RECT 2.080 0.318 2.141 0.486 ;
      RECT 2.040 0.318 2.080 0.475 ;
      RECT 1.953 0.171 2.043 0.252 ;
      RECT 1.743 0.420 2.040 0.475 ;
      RECT 1.926 0.198 1.953 0.252 ;
      RECT 1.845 0.795 1.936 0.876 ;
      RECT 1.865 0.198 1.926 0.325 ;
      RECT 1.493 0.270 1.865 0.325 ;
      RECT 1.743 0.795 1.845 0.850 ;
      RECT 1.682 0.420 1.743 0.850 ;
      RECT 1.579 0.426 1.682 0.507 ;
      RECT 1.560 0.563 1.621 0.917 ;
      RECT 1.491 0.563 1.560 0.618 ;
      RECT 1.425 0.862 1.560 0.917 ;
      RECT 1.409 0.700 1.499 0.781 ;
      RECT 1.491 0.204 1.493 0.325 ;
      RECT 1.430 0.204 1.491 0.618 ;
      RECT 1.409 0.204 1.430 0.271 ;
      RECT 1.335 0.862 1.425 0.943 ;
      RECT 1.319 0.190 1.409 0.271 ;
      RECT 1.326 0.700 1.409 0.755 ;
      RECT 1.326 0.438 1.340 0.519 ;
      RECT 1.265 0.438 1.326 0.755 ;
      RECT 1.250 0.438 1.265 0.519 ;
      RECT 0.978 0.601 1.265 0.656 ;
      RECT 1.123 0.825 1.213 0.906 ;
      RECT 1.183 0.257 1.196 0.338 ;
      RECT 1.106 0.206 1.183 0.338 ;
      RECT 0.863 0.851 1.123 0.906 ;
      RECT 0.457 0.206 1.106 0.261 ;
      RECT 0.917 0.601 0.978 0.787 ;
      RECT 0.740 0.732 0.917 0.787 ;
      RECT 0.802 0.851 0.863 1.025 ;
      RECT 0.438 0.970 0.802 1.025 ;
      RECT 0.679 0.732 0.740 0.915 ;
      RECT 0.138 0.861 0.679 0.915 ;
      RECT 0.557 0.389 0.618 0.789 ;
      RECT 0.536 0.389 0.557 0.444 ;
      RECT 0.404 0.735 0.557 0.789 ;
      RECT 0.460 0.346 0.536 0.444 ;
      RECT 0.445 0.346 0.460 0.427 ;
      RECT 0.396 0.152 0.457 0.261 ;
      RECT 0.098 0.331 0.138 0.412 ;
      RECT 0.098 0.743 0.138 0.915 ;
      RECT 0.077 0.331 0.098 0.915 ;
      RECT 0.048 0.331 0.077 0.824 ;
      RECT 0.037 0.331 0.048 0.807 ;
  END
END SDFFSHQX1

MACRO SDFFSXL
  CLASS CORE ;
  FOREIGN SDFFSXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.187 0.967 3.354 1.050 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.835 0.502 0.868 0.627 ;
      RECT 0.807 0.502 0.835 0.631 ;
      RECT 0.729 0.512 0.807 0.631 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.220 0.432 0.424 0.500 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.765 0.206 3.826 0.940 ;
      RECT 3.639 0.206 3.765 0.261 ;
      RECT 3.712 0.886 3.765 0.940 ;
      RECT 3.618 0.886 3.712 0.977 ;
      RECT 3.578 0.162 3.639 0.261 ;
      RECT 3.557 0.886 3.618 1.027 ;
      RECT 3.521 0.162 3.578 0.243 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.968 0.736 4.046 0.817 ;
      RECT 3.968 0.298 4.036 0.379 ;
      RECT 3.945 0.298 3.968 0.817 ;
      RECT 3.907 0.311 3.945 0.817 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.188 0.495 1.196 0.550 ;
      RECT 1.087 0.433 1.188 0.560 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.674 0.200 0.767 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.863 -0.080 4.200 0.080 ;
      RECT 3.773 -0.080 3.863 0.122 ;
      RECT 3.410 -0.080 3.773 0.080 ;
      RECT 3.320 -0.080 3.410 0.122 ;
      RECT 3.023 -0.080 3.320 0.080 ;
      RECT 2.933 -0.080 3.023 0.122 ;
      RECT 2.388 -0.080 2.933 0.080 ;
      RECT 2.327 -0.080 2.388 0.192 ;
      RECT 1.851 -0.080 2.327 0.080 ;
      RECT 1.761 -0.080 1.851 0.222 ;
      RECT 0.951 -0.080 1.761 0.080 ;
      RECT 0.860 -0.080 0.951 0.122 ;
      RECT 0.378 -0.080 0.860 0.080 ;
      RECT 0.288 -0.080 0.378 0.122 ;
      RECT 0.000 -0.080 0.288 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.910 1.120 4.200 1.280 ;
      RECT 3.804 1.078 3.910 1.280 ;
      RECT 3.476 1.120 3.804 1.280 ;
      RECT 3.476 0.710 3.521 0.761 ;
      RECT 3.431 0.710 3.476 1.280 ;
      RECT 3.415 0.723 3.431 1.280 ;
      RECT 3.126 1.120 3.415 1.280 ;
      RECT 3.036 1.001 3.126 1.280 ;
      RECT 2.461 1.120 3.036 1.280 ;
      RECT 2.370 1.001 2.461 1.280 ;
      RECT 2.112 1.120 2.370 1.280 ;
      RECT 2.051 1.001 2.112 1.280 ;
      RECT 1.755 1.120 2.051 1.280 ;
      RECT 1.665 1.078 1.755 1.280 ;
      RECT 0.924 1.120 1.665 1.280 ;
      RECT 0.863 0.991 0.924 1.280 ;
      RECT 0.286 1.120 0.863 1.280 ;
      RECT 0.196 1.078 0.286 1.280 ;
      RECT 0.000 1.120 0.196 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.698 0.368 3.704 0.700 ;
      RECT 3.643 0.368 3.698 0.776 ;
      RECT 3.622 0.368 3.643 0.423 ;
      RECT 3.637 0.645 3.643 0.776 ;
      RECT 3.532 0.342 3.622 0.423 ;
      RECT 3.320 0.482 3.541 0.537 ;
      RECT 3.268 0.451 3.320 0.805 ;
      RECT 3.259 0.361 3.268 0.805 ;
      RECT 3.207 0.361 3.259 0.506 ;
      RECT 3.230 0.724 3.259 0.805 ;
      RECT 3.102 0.361 3.207 0.415 ;
      RECT 2.796 0.580 3.192 0.635 ;
      RECT 3.012 0.335 3.102 0.415 ;
      RECT 2.930 0.335 3.012 0.389 ;
      RECT 2.868 0.276 2.930 0.389 ;
      RECT 2.840 0.276 2.868 0.357 ;
      RECT 2.796 0.783 2.811 0.864 ;
      RECT 2.777 0.446 2.796 0.864 ;
      RECT 2.735 0.356 2.777 0.864 ;
      RECT 2.718 0.356 2.735 0.501 ;
      RECT 2.720 0.783 2.735 0.864 ;
      RECT 2.716 0.343 2.718 0.501 ;
      RECT 2.628 0.343 2.716 0.424 ;
      RECT 2.622 0.957 2.713 1.038 ;
      RECT 2.592 0.480 2.636 0.561 ;
      RECT 2.583 0.957 2.622 1.012 ;
      RECT 2.567 0.480 2.592 0.749 ;
      RECT 2.522 0.874 2.583 1.012 ;
      RECT 2.506 0.296 2.567 0.749 ;
      RECT 1.656 0.874 2.522 0.929 ;
      RECT 2.266 0.296 2.506 0.351 ;
      RECT 2.313 0.694 2.506 0.749 ;
      RECT 2.353 0.515 2.443 0.596 ;
      RECT 2.191 0.529 2.353 0.583 ;
      RECT 2.252 0.694 2.313 0.814 ;
      RECT 2.205 0.173 2.266 0.351 ;
      RECT 2.130 0.173 2.205 0.227 ;
      RECT 2.144 0.529 2.191 0.813 ;
      RECT 2.130 0.345 2.144 0.813 ;
      RECT 2.070 0.151 2.130 0.227 ;
      RECT 2.083 0.345 2.130 0.583 ;
      RECT 1.716 0.758 2.130 0.813 ;
      RECT 1.938 0.151 2.070 0.206 ;
      RECT 1.917 0.582 2.007 0.663 ;
      RECT 1.838 0.582 1.917 0.637 ;
      RECT 1.777 0.519 1.838 0.637 ;
      RECT 1.509 0.519 1.777 0.574 ;
      RECT 1.655 0.629 1.716 0.813 ;
      RECT 1.595 0.874 1.656 0.973 ;
      RECT 1.623 0.629 1.655 0.683 ;
      RECT 1.507 0.918 1.595 0.973 ;
      RECT 1.509 0.162 1.523 0.243 ;
      RECT 1.448 0.162 1.509 0.744 ;
      RECT 1.432 0.918 1.507 1.049 ;
      RECT 1.433 0.162 1.448 0.243 ;
      RECT 1.444 0.689 1.448 0.744 ;
      RECT 1.383 0.689 1.444 0.838 ;
      RECT 1.322 0.994 1.432 1.049 ;
      RECT 1.371 0.333 1.385 0.414 ;
      RECT 1.322 0.333 1.371 0.579 ;
      RECT 1.310 0.333 1.322 1.049 ;
      RECT 1.221 0.181 1.311 0.262 ;
      RECT 1.295 0.333 1.310 0.414 ;
      RECT 1.261 0.524 1.310 1.049 ;
      RECT 1.046 0.994 1.261 1.049 ;
      RECT 0.700 0.207 1.221 0.262 ;
      RECT 1.168 0.885 1.200 0.939 ;
      RECT 1.107 0.723 1.168 0.939 ;
      RECT 0.643 0.723 1.107 0.777 ;
      RECT 0.985 0.864 1.046 1.049 ;
      RECT 0.640 0.335 1.025 0.389 ;
      RECT 0.801 0.864 0.985 0.919 ;
      RECT 0.740 0.864 0.801 1.039 ;
      RECT 0.447 0.985 0.740 1.039 ;
      RECT 0.639 0.165 0.700 0.262 ;
      RECT 0.640 0.587 0.655 0.668 ;
      RECT 0.631 0.723 0.643 0.915 ;
      RECT 0.590 0.335 0.640 0.668 ;
      RECT 0.500 0.165 0.639 0.220 ;
      RECT 0.582 0.723 0.631 0.929 ;
      RECT 0.579 0.321 0.590 0.668 ;
      RECT 0.541 0.848 0.582 0.929 ;
      RECT 0.500 0.321 0.579 0.402 ;
      RECT 0.565 0.587 0.579 0.668 ;
      RECT 0.484 0.613 0.565 0.668 ;
      RECT 0.423 0.613 0.484 0.752 ;
      RECT 0.386 0.869 0.447 1.039 ;
      RECT 0.322 0.869 0.386 0.924 ;
      RECT 0.261 0.560 0.322 0.924 ;
      RECT 0.109 0.560 0.261 0.614 ;
      RECT 0.048 0.843 0.261 0.924 ;
      RECT 0.109 0.283 0.138 0.364 ;
      RECT 0.048 0.283 0.109 0.614 ;
  END
END SDFFSXL

MACRO SDFFSX4
  CLASS CORE ;
  FOREIGN SDFFSX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.901 0.962 2.063 1.050 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.756 0.488 0.862 0.627 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.433 0.468 0.595 ;
      RECT 0.374 0.494 0.387 0.595 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.038 0.324 5.043 0.405 ;
      RECT 5.038 0.652 5.043 0.733 ;
      RECT 4.948 0.300 5.038 0.733 ;
      RECT 4.937 0.300 4.948 0.633 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.523 0.433 5.563 0.767 ;
      RECT 5.462 0.350 5.523 0.767 ;
      RECT 5.383 0.350 5.462 0.405 ;
      RECT 5.292 0.652 5.462 0.733 ;
      RECT 5.292 0.324 5.383 0.405 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.054 0.438 1.168 0.563 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.252 0.567 0.313 0.633 ;
      RECT 0.191 0.437 0.252 0.633 ;
      RECT 0.162 0.437 0.191 0.518 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.552 -0.080 5.600 0.080 ;
      RECT 5.462 -0.080 5.552 0.211 ;
      RECT 5.213 -0.080 5.462 0.080 ;
      RECT 5.123 -0.080 5.213 0.211 ;
      RECT 4.863 -0.080 5.123 0.080 ;
      RECT 4.773 -0.080 4.863 0.122 ;
      RECT 4.505 -0.080 4.773 0.080 ;
      RECT 4.415 -0.080 4.505 0.247 ;
      RECT 3.816 -0.080 4.415 0.080 ;
      RECT 3.725 -0.080 3.816 0.122 ;
      RECT 3.288 -0.080 3.725 0.080 ;
      RECT 3.198 -0.080 3.288 0.299 ;
      RECT 2.609 -0.080 3.198 0.080 ;
      RECT 2.519 -0.080 2.609 0.299 ;
      RECT 1.835 -0.080 2.519 0.080 ;
      RECT 1.745 -0.080 1.835 0.290 ;
      RECT 0.902 -0.080 1.745 0.080 ;
      RECT 0.811 -0.080 0.902 0.122 ;
      RECT 0.313 -0.080 0.811 0.080 ;
      RECT 0.223 -0.080 0.313 0.122 ;
      RECT 0.000 -0.080 0.223 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.552 1.120 5.600 1.280 ;
      RECT 5.462 0.989 5.552 1.280 ;
      RECT 5.213 1.120 5.462 1.280 ;
      RECT 5.123 0.989 5.213 1.280 ;
      RECT 4.863 1.120 5.123 1.280 ;
      RECT 4.773 1.078 4.863 1.280 ;
      RECT 4.484 1.120 4.773 1.280 ;
      RECT 4.394 0.779 4.484 1.280 ;
      RECT 4.102 1.120 4.394 1.280 ;
      RECT 4.012 0.833 4.102 1.280 ;
      RECT 3.709 1.120 4.012 1.280 ;
      RECT 3.619 0.977 3.709 1.280 ;
      RECT 3.256 1.120 3.619 1.280 ;
      RECT 3.166 0.971 3.256 1.280 ;
      RECT 2.556 1.120 3.166 1.280 ;
      RECT 2.466 0.971 2.556 1.280 ;
      RECT 2.186 1.120 2.466 1.280 ;
      RECT 2.125 0.971 2.186 1.280 ;
      RECT 1.836 1.120 2.125 1.280 ;
      RECT 1.775 1.003 1.836 1.280 ;
      RECT 0.941 1.120 1.775 1.280 ;
      RECT 0.851 1.001 0.941 1.280 ;
      RECT 0.198 1.120 0.851 1.280 ;
      RECT 0.065 1.077 0.198 1.280 ;
      RECT 0.000 1.120 0.065 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.220 0.486 5.284 0.567 ;
      RECT 5.194 0.486 5.220 0.888 ;
      RECT 5.159 0.512 5.194 0.888 ;
      RECT 4.696 0.833 5.159 0.888 ;
      RECT 4.635 0.305 4.696 0.888 ;
      RECT 4.606 0.305 4.635 0.386 ;
      RECT 4.584 0.807 4.635 0.888 ;
      RECT 4.484 0.495 4.574 0.576 ;
      RECT 4.293 0.496 4.484 0.575 ;
      RECT 4.232 0.358 4.293 0.845 ;
      RECT 4.166 0.358 4.232 0.413 ;
      RECT 4.203 0.708 4.232 0.845 ;
      RECT 3.911 0.708 4.203 0.763 ;
      RECT 4.109 0.295 4.166 0.413 ;
      RECT 4.048 0.251 4.109 0.413 ;
      RECT 4.012 0.507 4.102 0.588 ;
      RECT 3.638 0.251 4.048 0.306 ;
      RECT 3.476 0.520 4.012 0.575 ;
      RECT 3.850 0.708 3.911 0.887 ;
      RECT 3.821 0.768 3.850 0.887 ;
      RECT 3.538 0.832 3.821 0.887 ;
      RECT 3.477 0.832 3.538 0.963 ;
      RECT 3.415 0.340 3.476 0.745 ;
      RECT 3.386 0.340 3.415 0.424 ;
      RECT 3.402 0.690 3.415 0.745 ;
      RECT 3.312 0.690 3.402 0.771 ;
      RECT 3.135 0.369 3.386 0.424 ;
      RECT 3.253 0.529 3.344 0.610 ;
      RECT 2.906 0.704 3.312 0.758 ;
      RECT 2.999 0.542 3.253 0.596 ;
      RECT 3.074 0.270 3.135 0.424 ;
      RECT 2.948 0.270 3.074 0.325 ;
      RECT 2.938 0.407 2.999 0.596 ;
      RECT 2.858 0.257 2.948 0.338 ;
      RECT 2.909 0.407 2.938 0.488 ;
      RECT 2.595 0.420 2.909 0.475 ;
      RECT 2.816 0.704 2.906 0.819 ;
      RECT 2.732 0.530 2.821 0.585 ;
      RECT 2.671 0.530 2.732 0.901 ;
      RECT 2.349 0.846 2.671 0.901 ;
      RECT 2.534 0.420 2.595 0.777 ;
      RECT 2.397 0.420 2.534 0.475 ;
      RECT 2.402 0.723 2.534 0.777 ;
      RECT 2.378 0.540 2.469 0.621 ;
      RECT 2.312 0.710 2.402 0.790 ;
      RECT 2.356 0.276 2.397 0.475 ;
      RECT 2.221 0.554 2.378 0.608 ;
      RECT 2.321 0.150 2.356 0.475 ;
      RECT 2.259 0.846 2.349 0.955 ;
      RECT 2.295 0.150 2.321 0.357 ;
      RECT 2.282 0.150 2.295 0.231 ;
      RECT 1.645 0.846 2.259 0.901 ;
      RECT 2.174 0.273 2.221 0.764 ;
      RECT 2.160 0.229 2.174 0.764 ;
      RECT 2.084 0.229 2.160 0.327 ;
      RECT 2.052 0.710 2.160 0.764 ;
      RECT 1.986 0.382 2.076 0.463 ;
      RECT 1.962 0.710 2.052 0.790 ;
      RECT 1.525 0.382 1.986 0.437 ;
      RECT 1.847 0.710 1.962 0.764 ;
      RECT 1.786 0.518 1.847 0.764 ;
      RECT 1.761 0.518 1.786 0.573 ;
      RECT 1.670 0.492 1.761 0.573 ;
      RECT 1.584 0.846 1.645 1.020 ;
      RECT 1.401 0.965 1.584 1.020 ;
      RECT 1.523 0.261 1.525 0.437 ;
      RECT 1.474 0.261 1.523 0.886 ;
      RECT 1.462 0.248 1.474 0.886 ;
      RECT 1.384 0.248 1.462 0.329 ;
      RECT 1.400 0.396 1.401 1.020 ;
      RECT 1.340 0.383 1.400 1.020 ;
      RECT 1.310 0.383 1.340 0.464 ;
      RECT 1.156 0.693 1.340 0.748 ;
      RECT 1.218 0.805 1.279 0.931 ;
      RECT 1.172 0.185 1.262 0.265 ;
      RECT 0.790 0.876 1.218 0.931 ;
      RECT 0.705 0.205 1.172 0.260 ;
      RECT 1.095 0.693 1.156 0.821 ;
      RECT 0.668 0.767 1.095 0.821 ;
      RECT 0.640 0.324 0.976 0.379 ;
      RECT 0.729 0.876 0.790 0.958 ;
      RECT 0.491 0.904 0.729 0.958 ;
      RECT 0.644 0.155 0.705 0.260 ;
      RECT 0.607 0.767 0.668 0.849 ;
      RECT 0.640 0.631 0.655 0.712 ;
      RECT 0.451 0.155 0.644 0.210 ;
      RECT 0.579 0.324 0.640 0.712 ;
      RECT 0.159 0.794 0.607 0.849 ;
      RECT 0.435 0.324 0.579 0.379 ;
      RECT 0.565 0.631 0.579 0.712 ;
      RECT 0.514 0.657 0.565 0.712 ;
      RECT 0.424 0.657 0.514 0.739 ;
      RECT 0.101 0.299 0.159 0.380 ;
      RECT 0.101 0.705 0.159 0.849 ;
      RECT 0.098 0.299 0.101 0.849 ;
      RECT 0.040 0.299 0.098 0.786 ;
  END
END SDFFSX4

MACRO SDFFRHQXL
  CLASS CORE ;
  FOREIGN SDFFRHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.877 0.567 0.999 0.627 ;
      RECT 0.801 0.488 0.877 0.627 ;
      RECT 0.787 0.488 0.801 0.569 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.380 0.433 0.499 0.543 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.987 0.706 3.991 0.761 ;
      RECT 3.776 0.693 3.987 0.776 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.363 0.302 4.367 0.761 ;
      RECT 4.305 0.302 4.363 0.965 ;
      RECT 4.077 0.302 4.305 0.357 ;
      RECT 4.281 0.706 4.305 0.965 ;
      RECT 4.256 0.885 4.281 0.965 ;
      RECT 4.016 0.167 4.077 0.357 ;
      RECT 3.987 0.167 4.016 0.248 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.035 0.417 1.195 0.502 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.233 0.517 0.295 0.627 ;
      RECT 0.168 0.517 0.233 0.625 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.291 -0.080 4.400 0.080 ;
      RECT 4.200 -0.080 4.291 0.233 ;
      RECT 3.863 -0.080 4.200 0.080 ;
      RECT 3.612 -0.080 3.863 0.122 ;
      RECT 3.308 -0.080 3.612 0.080 ;
      RECT 3.217 -0.080 3.308 0.122 ;
      RECT 2.515 -0.080 3.217 0.080 ;
      RECT 2.424 -0.080 2.515 0.261 ;
      RECT 1.797 -0.080 2.424 0.080 ;
      RECT 2.144 0.363 2.173 0.414 ;
      RECT 2.083 0.288 2.144 0.414 ;
      RECT 1.797 0.288 2.083 0.338 ;
      RECT 1.707 -0.080 1.797 0.338 ;
      RECT 0.868 -0.080 1.707 0.080 ;
      RECT 0.777 -0.080 0.868 0.122 ;
      RECT 0.301 -0.080 0.777 0.080 ;
      RECT 0.211 -0.080 0.301 0.122 ;
      RECT 0.000 -0.080 0.211 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.005 1.120 4.400 1.280 ;
      RECT 3.915 0.850 4.005 1.280 ;
      RECT 3.395 1.120 3.915 1.280 ;
      RECT 3.284 1.078 3.395 1.280 ;
      RECT 2.605 1.120 3.284 1.280 ;
      RECT 2.515 1.078 2.605 1.280 ;
      RECT 1.781 1.120 2.515 1.280 ;
      RECT 1.691 0.967 1.781 1.280 ;
      RECT 0.933 1.120 1.691 1.280 ;
      RECT 0.843 0.998 0.933 1.280 ;
      RECT 0.245 1.120 0.843 1.280 ;
      RECT 0.155 0.928 0.245 1.280 ;
      RECT 0.000 1.120 0.155 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.851 0.420 4.219 0.475 ;
      RECT 3.681 0.581 4.068 0.636 ;
      RECT 3.789 0.206 3.851 0.475 ;
      RECT 3.537 0.944 3.792 0.999 ;
      RECT 3.404 0.206 3.789 0.261 ;
      RECT 3.681 0.327 3.703 0.408 ;
      RECT 3.673 0.327 3.681 0.636 ;
      RECT 3.612 0.327 3.673 0.638 ;
      RECT 3.537 0.526 3.612 0.638 ;
      RECT 3.527 0.526 3.537 0.999 ;
      RECT 3.476 0.573 3.527 0.999 ;
      RECT 3.399 0.336 3.489 0.417 ;
      RECT 2.247 0.944 3.476 0.999 ;
      RECT 3.305 0.206 3.404 0.273 ;
      RECT 3.381 0.362 3.399 0.417 ;
      RECT 3.320 0.362 3.381 0.820 ;
      RECT 3.269 0.605 3.320 0.820 ;
      RECT 3.164 0.206 3.305 0.261 ;
      RECT 3.225 0.605 3.269 0.688 ;
      RECT 3.103 0.206 3.164 0.857 ;
      RECT 2.944 0.206 3.103 0.263 ;
      RECT 3.016 0.802 3.103 0.857 ;
      RECT 2.965 0.383 3.019 0.464 ;
      RECT 2.925 0.802 3.016 0.883 ;
      RECT 2.904 0.383 2.965 0.727 ;
      RECT 2.853 0.206 2.944 0.306 ;
      RECT 2.824 0.380 2.843 0.870 ;
      RECT 2.788 0.380 2.824 0.883 ;
      RECT 2.781 0.249 2.788 0.883 ;
      RECT 2.731 0.249 2.781 0.435 ;
      RECT 2.733 0.802 2.781 0.883 ;
      RECT 2.727 0.236 2.731 0.435 ;
      RECT 2.640 0.236 2.727 0.317 ;
      RECT 2.660 0.543 2.720 0.624 ;
      RECT 2.599 0.388 2.660 0.829 ;
      RECT 2.403 0.388 2.599 0.443 ;
      RECT 2.472 0.774 2.599 0.829 ;
      RECT 2.508 0.613 2.537 0.694 ;
      RECT 2.447 0.525 2.508 0.694 ;
      RECT 2.381 0.774 2.472 0.855 ;
      RECT 2.001 0.525 2.447 0.580 ;
      RECT 2.359 0.362 2.403 0.443 ;
      RECT 2.297 0.163 2.359 0.443 ;
      RECT 1.867 0.163 2.297 0.218 ;
      RECT 2.185 0.638 2.247 0.999 ;
      RECT 2.123 0.638 2.185 0.719 ;
      RECT 1.940 0.389 2.001 0.876 ;
      RECT 1.689 0.389 1.940 0.451 ;
      RECT 1.880 0.795 1.940 0.876 ;
      RECT 1.788 0.627 1.879 0.711 ;
      RECT 1.487 0.656 1.788 0.711 ;
      RECT 1.628 0.389 1.689 0.564 ;
      RECT 1.599 0.483 1.628 0.564 ;
      RECT 1.459 0.890 1.549 0.971 ;
      RECT 1.449 0.226 1.487 0.711 ;
      RECT 1.319 0.890 1.459 0.945 ;
      RECT 1.425 0.226 1.449 0.792 ;
      RECT 1.424 0.226 1.425 0.281 ;
      RECT 1.388 0.646 1.425 0.792 ;
      RECT 1.333 0.200 1.424 0.281 ;
      RECT 1.257 0.394 1.319 0.945 ;
      RECT 0.629 0.732 1.257 0.787 ;
      RECT 1.141 0.195 1.232 0.276 ;
      RECT 1.135 0.856 1.196 0.996 ;
      RECT 0.508 0.208 1.141 0.263 ;
      RECT 0.756 0.856 1.135 0.911 ;
      RECT 0.853 0.327 0.944 0.408 ;
      RECT 0.629 0.354 0.853 0.408 ;
      RECT 0.695 0.856 0.756 0.967 ;
      RECT 0.533 0.912 0.695 0.967 ;
      RECT 0.629 0.595 0.691 0.676 ;
      RECT 0.568 0.348 0.629 0.676 ;
      RECT 0.568 0.732 0.629 0.857 ;
      RECT 0.491 0.621 0.568 0.676 ;
      RECT 0.324 0.802 0.568 0.857 ;
      RECT 0.447 0.150 0.508 0.263 ;
      RECT 0.429 0.621 0.491 0.748 ;
      RECT 0.397 0.150 0.447 0.205 ;
      RECT 0.400 0.667 0.429 0.748 ;
      RECT 0.263 0.688 0.324 0.857 ;
      RECT 0.139 0.688 0.263 0.743 ;
      RECT 0.105 0.333 0.139 0.414 ;
      RECT 0.105 0.680 0.139 0.743 ;
      RECT 0.044 0.333 0.105 0.743 ;
  END
END SDFFRHQXL

MACRO SDFFRHQX4
  CLASS CORE ;
  FOREIGN SDFFRHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.729 0.671 0.828 0.806 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.981 0.562 1.090 0.617 ;
      RECT 0.921 0.562 0.981 0.627 ;
      RECT 0.829 0.562 0.921 0.617 ;
      RECT 0.769 0.454 0.829 0.617 ;
      RECT 0.689 0.454 0.769 0.508 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.529 0.437 4.787 0.500 ;
      RECT 4.527 0.437 4.529 0.492 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 6.319 0.707 6.333 0.931 ;
      RECT 6.244 0.706 6.319 0.931 ;
      RECT 6.190 0.706 6.244 0.767 ;
      RECT 6.091 0.349 6.190 0.767 ;
      RECT 6.007 0.349 6.091 0.404 ;
      RECT 5.662 0.712 6.091 0.767 ;
      RECT 5.918 0.179 6.007 0.404 ;
      RECT 5.629 0.349 5.918 0.404 ;
      RECT 5.573 0.707 5.662 0.931 ;
      RECT 5.555 0.179 5.629 0.404 ;
      RECT 5.540 0.179 5.555 0.402 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 0.706 1.206 0.792 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.165 0.476 0.290 0.627 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.196 -0.080 6.400 0.080 ;
      RECT 6.106 -0.080 6.196 0.235 ;
      RECT 5.818 -0.080 6.106 0.080 ;
      RECT 5.729 -0.080 5.818 0.235 ;
      RECT 5.377 -0.080 5.729 0.080 ;
      RECT 5.316 -0.080 5.377 0.360 ;
      RECT 4.923 -0.080 5.316 0.080 ;
      RECT 4.834 -0.080 4.923 0.122 ;
      RECT 4.535 -0.080 4.834 0.080 ;
      RECT 4.446 -0.080 4.535 0.268 ;
      RECT 3.083 -0.080 4.446 0.080 ;
      RECT 2.994 -0.080 3.083 0.299 ;
      RECT 2.706 -0.080 2.994 0.080 ;
      RECT 2.617 -0.080 2.706 0.340 ;
      RECT 2.267 -0.080 2.617 0.080 ;
      RECT 2.267 0.315 2.281 0.366 ;
      RECT 2.207 -0.080 2.267 0.366 ;
      RECT 1.894 -0.080 2.207 0.080 ;
      RECT 2.192 0.315 2.207 0.366 ;
      RECT 1.804 -0.080 1.894 0.216 ;
      RECT 1.051 -0.080 1.804 0.080 ;
      RECT 0.962 -0.080 1.051 0.122 ;
      RECT 0.337 -0.080 0.962 0.080 ;
      RECT 0.248 -0.080 0.337 0.122 ;
      RECT 0.000 -0.080 0.248 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.998 1.120 6.400 1.280 ;
      RECT 5.909 0.910 5.998 1.280 ;
      RECT 5.312 1.120 5.909 1.280 ;
      RECT 5.252 0.742 5.312 1.280 ;
      RECT 4.881 1.120 5.252 1.280 ;
      RECT 4.792 1.078 4.881 1.280 ;
      RECT 4.450 1.120 4.792 1.280 ;
      RECT 4.361 0.989 4.450 1.280 ;
      RECT 3.141 1.120 4.361 1.280 ;
      RECT 3.052 1.078 3.141 1.280 ;
      RECT 2.741 1.120 3.052 1.280 ;
      RECT 2.681 0.982 2.741 1.280 ;
      RECT 2.368 1.120 2.681 1.280 ;
      RECT 2.279 1.078 2.368 1.280 ;
      RECT 1.873 1.120 2.279 1.280 ;
      RECT 1.783 1.078 1.873 1.280 ;
      RECT 0.346 1.120 1.783 1.280 ;
      RECT 0.257 1.078 0.346 1.280 ;
      RECT 0.000 1.120 0.257 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.314 0.506 5.902 0.561 ;
      RECT 5.256 0.506 5.314 0.594 ;
      RECT 5.196 0.192 5.256 0.594 ;
      RECT 4.724 0.192 5.196 0.246 ;
      RECT 5.192 0.539 5.196 0.594 ;
      RECT 5.132 0.539 5.192 0.994 ;
      RECT 5.075 0.301 5.135 0.423 ;
      RECT 4.573 0.939 5.132 0.994 ;
      RECT 4.944 0.368 5.075 0.423 ;
      RECT 5.011 0.524 5.071 0.885 ;
      RECT 4.707 0.830 5.011 0.885 ;
      RECT 4.884 0.368 4.944 0.775 ;
      RECT 4.467 0.611 4.884 0.665 ;
      RECT 4.649 0.192 4.724 0.317 ;
      RECT 4.647 0.751 4.707 0.885 ;
      RECT 4.635 0.236 4.649 0.317 ;
      RECT 4.345 0.751 4.647 0.806 ;
      RECT 4.513 0.862 4.573 0.994 ;
      RECT 4.292 0.862 4.513 0.917 ;
      RECT 4.407 0.524 4.467 0.665 ;
      RECT 4.252 0.524 4.407 0.579 ;
      RECT 4.285 0.649 4.345 0.806 ;
      RECT 4.231 0.862 4.292 1.039 ;
      RECT 4.143 0.649 4.285 0.704 ;
      RECT 3.262 0.985 4.231 1.039 ;
      RECT 4.143 0.262 4.179 0.343 ;
      RECT 4.111 0.762 4.171 0.915 ;
      RECT 4.083 0.161 4.143 0.704 ;
      RECT 3.414 0.861 4.111 0.915 ;
      RECT 3.801 0.161 4.083 0.215 ;
      RECT 4.010 0.627 4.083 0.704 ;
      RECT 3.686 0.627 4.010 0.682 ;
      RECT 3.923 0.285 3.990 0.339 ;
      RECT 3.863 0.285 3.923 0.458 ;
      RECT 3.549 0.737 3.900 0.792 ;
      RECT 3.613 0.404 3.863 0.458 ;
      RECT 3.712 0.161 3.801 0.329 ;
      RECT 3.324 0.161 3.712 0.215 ;
      RECT 3.626 0.600 3.686 0.682 ;
      RECT 3.549 0.285 3.613 0.458 ;
      RECT 3.488 0.285 3.549 0.792 ;
      RECT 3.469 0.285 3.488 0.458 ;
      RECT 3.474 0.692 3.488 0.792 ;
      RECT 3.117 0.692 3.474 0.746 ;
      RECT 3.258 0.285 3.469 0.339 ;
      RECT 3.353 0.815 3.414 0.915 ;
      RECT 3.336 0.421 3.397 0.580 ;
      RECT 2.982 0.815 3.353 0.870 ;
      RECT 2.982 0.525 3.336 0.580 ;
      RECT 3.201 0.954 3.262 1.039 ;
      RECT 3.197 0.285 3.258 0.425 ;
      RECT 2.862 0.954 3.201 1.008 ;
      RECT 2.895 0.370 3.197 0.425 ;
      RECT 3.057 0.660 3.117 0.746 ;
      RECT 2.922 0.525 2.982 0.870 ;
      RECT 2.724 0.525 2.922 0.580 ;
      RECT 2.834 0.270 2.895 0.425 ;
      RECT 2.802 0.808 2.862 1.008 ;
      RECT 2.806 0.270 2.834 0.351 ;
      RECT 2.564 0.808 2.802 0.863 ;
      RECT 2.724 0.655 2.739 0.736 ;
      RECT 2.664 0.423 2.724 0.736 ;
      RECT 2.516 0.423 2.664 0.477 ;
      RECT 2.650 0.655 2.664 0.736 ;
      RECT 2.542 0.919 2.602 1.005 ;
      RECT 2.504 0.546 2.564 0.863 ;
      RECT 2.308 0.919 2.542 0.974 ;
      RECT 2.487 0.300 2.516 0.477 ;
      RECT 2.177 0.546 2.504 0.601 ;
      RECT 2.456 0.161 2.487 0.477 ;
      RECT 2.427 0.161 2.456 0.381 ;
      RECT 2.116 0.699 2.443 0.792 ;
      RECT 2.331 0.161 2.427 0.215 ;
      RECT 2.247 0.919 2.308 0.994 ;
      RECT 1.624 0.939 2.247 0.994 ;
      RECT 2.056 0.294 2.116 0.792 ;
      RECT 2.018 0.294 2.056 0.381 ;
      RECT 2.053 0.698 2.056 0.792 ;
      RECT 1.924 0.698 2.053 0.779 ;
      RECT 1.900 0.480 1.993 0.615 ;
      RECT 1.815 0.698 1.924 0.752 ;
      RECT 1.616 0.480 1.900 0.535 ;
      RECT 1.755 0.612 1.815 0.752 ;
      RECT 1.726 0.612 1.755 0.693 ;
      RECT 1.624 0.650 1.638 0.731 ;
      RECT 1.563 0.650 1.624 0.994 ;
      RECT 1.572 0.480 1.616 0.563 ;
      RECT 1.572 0.214 1.587 0.295 ;
      RECT 1.512 0.214 1.572 0.563 ;
      RECT 1.549 0.650 1.563 0.731 ;
      RECT 1.326 0.874 1.563 0.932 ;
      RECT 1.498 0.214 1.512 0.295 ;
      RECT 1.485 0.508 1.512 0.563 ;
      RECT 1.424 0.508 1.485 0.818 ;
      RECT 1.386 0.350 1.447 0.437 ;
      RECT 1.309 0.208 1.401 0.275 ;
      RECT 1.326 0.382 1.386 0.437 ;
      RECT 1.266 0.382 1.326 0.932 ;
      RECT 0.695 0.208 1.309 0.263 ;
      RECT 0.545 0.987 1.300 1.042 ;
      RECT 0.667 0.877 1.266 0.932 ;
      RECT 1.001 0.344 1.090 0.431 ;
      RECT 0.529 0.344 1.001 0.399 ;
      RECT 0.605 0.208 0.695 0.287 ;
      RECT 0.607 0.775 0.667 0.932 ;
      RECT 0.136 0.775 0.607 0.830 ;
      RECT 0.485 0.885 0.545 1.042 ;
      RECT 0.529 0.476 0.544 0.557 ;
      RECT 0.469 0.256 0.529 0.720 ;
      RECT 0.451 0.885 0.485 0.939 ;
      RECT 0.422 0.256 0.469 0.311 ;
      RECT 0.455 0.476 0.469 0.557 ;
      RECT 0.440 0.665 0.469 0.720 ;
      RECT 0.104 0.167 0.136 0.360 ;
      RECT 0.104 0.729 0.136 0.952 ;
      RECT 0.043 0.167 0.104 0.952 ;
  END
END SDFFRHQX4

MACRO SDFFRHQX2
  CLASS CORE ;
  FOREIGN SDFFRHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.865 0.567 0.984 0.629 ;
      RECT 0.776 0.548 0.865 0.629 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.383 0.415 0.491 0.543 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.216 0.632 4.357 0.763 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.937 0.275 4.998 0.729 ;
      RECT 4.643 0.275 4.937 0.330 ;
      RECT 4.817 0.674 4.937 0.729 ;
      RECT 4.727 0.674 4.817 0.960 ;
      RECT 4.641 0.225 4.643 0.330 ;
      RECT 4.551 0.151 4.641 0.344 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.019 0.418 1.177 0.510 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.290 0.506 0.310 0.617 ;
      RECT 0.230 0.506 0.290 0.627 ;
      RECT 0.158 0.506 0.230 0.617 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.840 -0.080 5.200 0.080 ;
      RECT 4.751 -0.080 4.840 0.122 ;
      RECT 4.382 -0.080 4.751 0.080 ;
      RECT 4.135 -0.080 4.382 0.122 ;
      RECT 3.782 -0.080 4.135 0.080 ;
      RECT 3.693 -0.080 3.782 0.122 ;
      RECT 2.754 -0.080 3.693 0.080 ;
      RECT 2.664 -0.080 2.754 0.292 ;
      RECT 1.731 -0.080 2.664 0.080 ;
#      RECT 2.035 0.303 2.125 0.359 ;
#      RECT 1.731 0.303 2.035 0.353 ;
      RECT 1.670 -0.080 1.731 0.328 ;
      RECT 1.641 -0.080 1.670 0.327 ;
      RECT 0.826 -0.080 1.641 0.080 ;
      RECT 0.737 -0.080 0.826 0.122 ;
      RECT 0.284 -0.080 0.737 0.080 ;
      RECT 0.194 -0.080 0.284 0.122 ;
      RECT 0.000 -0.080 0.194 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 1.120 5.200 1.280 ;
      RECT 5.063 0.800 5.153 1.280 ;
      RECT 4.457 1.120 5.063 1.280 ;
      RECT 4.367 1.078 4.457 1.280 ;
      RECT 4.089 1.120 4.367 1.280 ;
      RECT 4.000 1.078 4.089 1.280 ;
      RECT 3.778 1.120 4.000 1.280 ;
      RECT 3.662 1.078 3.778 1.280 ;
      RECT 2.759 1.120 3.662 1.280 ;
      RECT 2.670 1.078 2.759 1.280 ;
      RECT 1.754 1.120 2.670 1.280 ;
      RECT 1.665 0.997 1.754 1.280 ;
      RECT 0.919 1.120 1.665 1.280 ;
      RECT 0.830 1.001 0.919 1.280 ;
      RECT 0.347 1.120 0.830 1.280 ;
      RECT 0.336 1.013 0.347 1.280 ;
      RECT 0.247 0.972 0.336 1.280 ;
      RECT 0.236 1.013 0.247 1.280 ;
      RECT 0.000 1.120 0.236 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.725 0.538 4.877 0.619 ;
      RECT 4.664 0.399 4.725 0.619 ;
      RECT 4.411 0.399 4.664 0.454 ;
      RECT 4.473 0.523 4.562 0.612 ;
      RECT 4.289 0.523 4.473 0.577 ;
      RECT 4.350 0.206 4.411 0.454 ;
      RECT 3.925 0.206 4.350 0.261 ;
      RECT 4.226 0.838 4.315 0.919 ;
      RECT 4.199 0.352 4.289 0.577 ;
      RECT 4.025 0.838 4.226 0.893 ;
      RECT 4.094 0.523 4.199 0.577 ;
      RECT 4.025 0.517 4.094 0.598 ;
      RECT 4.005 0.517 4.025 0.994 ;
      RECT 3.921 0.336 4.010 0.417 ;
      RECT 3.964 0.543 4.005 0.994 ;
      RECT 3.431 0.939 3.964 0.994 ;
      RECT 3.832 0.206 3.925 0.273 ;
      RECT 3.807 0.349 3.921 0.404 ;
      RECT 3.425 0.206 3.832 0.261 ;
      RECT 3.807 0.736 3.821 0.817 ;
      RECT 3.746 0.349 3.807 0.817 ;
      RECT 3.732 0.605 3.746 0.817 ;
      RECT 3.658 0.605 3.732 0.686 ;
      RECT 3.484 0.360 3.498 0.440 ;
      RECT 3.459 0.360 3.484 0.688 ;
      RECT 3.423 0.360 3.459 0.714 ;
      RECT 3.371 0.939 3.431 1.039 ;
      RECT 3.334 0.170 3.425 0.261 ;
      RECT 3.409 0.360 3.423 0.440 ;
      RECT 3.369 0.633 3.423 0.714 ;
      RECT 2.916 0.985 3.371 1.039 ;
      RECT 3.310 0.795 3.362 0.876 ;
      RECT 3.158 0.206 3.334 0.261 ;
      RECT 3.305 0.338 3.325 0.419 ;
      RECT 3.305 0.795 3.310 0.915 ;
      RECT 3.245 0.338 3.305 0.915 ;
      RECT 3.236 0.338 3.245 0.419 ;
      RECT 3.037 0.861 3.245 0.915 ;
      RECT 3.098 0.206 3.158 0.786 ;
      RECT 3.058 0.206 3.098 0.419 ;
      RECT 2.983 0.817 3.037 0.915 ;
      RECT 2.977 0.804 2.983 0.915 ;
      RECT 2.968 0.804 2.977 0.885 ;
      RECT 2.943 0.362 2.968 0.885 ;
      RECT 2.907 0.240 2.943 0.885 ;
      RECT 2.856 0.939 2.916 1.039 ;
      RECT 2.853 0.240 2.907 0.417 ;
      RECT 2.894 0.804 2.907 0.885 ;
      RECT 2.621 0.817 2.894 0.871 ;
      RECT 2.184 0.939 2.856 0.994 ;
      RECT 2.550 0.362 2.853 0.417 ;
      RECT 2.786 0.471 2.847 0.746 ;
      RECT 2.428 0.471 2.786 0.526 ;
      RECT 2.437 0.692 2.786 0.746 ;
      RECT 2.307 0.582 2.684 0.637 ;
      RECT 2.532 0.802 2.621 0.883 ;
      RECT 2.490 0.252 2.550 0.417 ;
      RECT 2.377 0.692 2.437 0.829 ;
      RECT 2.368 0.319 2.428 0.526 ;
      RECT 2.348 0.748 2.377 0.829 ;
      RECT 2.336 0.319 2.368 0.374 ;
      RECT 2.307 0.293 2.336 0.374 ;
      RECT 2.247 0.176 2.307 0.374 ;
      RECT 2.247 0.477 2.307 0.637 ;
      RECT 1.901 0.176 2.247 0.231 ;
      RECT 1.976 0.477 2.247 0.532 ;
      RECT 2.123 0.607 2.184 0.994 ;
      RECT 1.916 0.477 1.976 0.876 ;
      RECT 1.915 0.477 1.916 0.532 ;
      RECT 1.853 0.795 1.916 0.876 ;
      RECT 1.825 0.398 1.915 0.532 ;
      RECT 1.812 0.150 1.901 0.231 ;
      RECT 1.743 0.607 1.832 0.701 ;
      RECT 1.656 0.477 1.825 0.532 ;
      RECT 1.454 0.646 1.743 0.701 ;
      RECT 1.595 0.477 1.656 0.590 ;
      RECT 1.567 0.510 1.595 0.590 ;
      RECT 1.494 0.902 1.509 0.983 ;
      RECT 1.419 0.901 1.494 0.983 ;
      RECT 1.393 0.176 1.454 0.792 ;
      RECT 1.299 0.901 1.419 0.956 ;
      RECT 1.372 0.176 1.393 0.231 ;
      RECT 1.359 0.698 1.393 0.792 ;
      RECT 1.283 0.150 1.372 0.231 ;
      RECT 1.299 0.445 1.301 0.630 ;
      RECT 1.241 0.445 1.299 0.956 ;
      RECT 1.238 0.575 1.241 0.956 ;
      RECT 0.599 0.732 1.238 0.787 ;
      RECT 1.098 0.202 1.187 0.283 ;
      RECT 1.117 0.856 1.178 0.995 ;
      RECT 0.755 0.856 1.117 0.911 ;
      RECT 0.545 0.206 1.098 0.261 ;
      RECT 0.852 0.324 0.901 0.405 ;
      RECT 0.624 0.323 0.852 0.405 ;
      RECT 0.695 0.856 0.755 0.993 ;
      RECT 0.615 0.938 0.695 0.993 ;
      RECT 0.624 0.595 0.688 0.676 ;
      RECT 0.599 0.323 0.624 0.676 ;
      RECT 0.525 0.938 0.615 1.019 ;
      RECT 0.552 0.323 0.599 0.663 ;
      RECT 0.538 0.732 0.599 0.858 ;
      RECT 0.469 0.608 0.552 0.663 ;
      RECT 0.485 0.165 0.545 0.261 ;
      RECT 0.137 0.804 0.538 0.858 ;
      RECT 0.378 0.165 0.485 0.220 ;
      RECT 0.408 0.608 0.469 0.748 ;
      RECT 0.122 0.318 0.137 0.399 ;
      RECT 0.097 0.671 0.137 0.864 ;
      RECT 0.097 0.318 0.122 0.450 ;
      RECT 0.047 0.318 0.097 0.864 ;
      RECT 0.037 0.395 0.047 0.726 ;
  END
END SDFFRHQX2

MACRO SDFFRHQX1
  CLASS CORE ;
  FOREIGN SDFFRHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.877 0.567 0.999 0.627 ;
      RECT 0.801 0.488 0.877 0.627 ;
      RECT 0.787 0.488 0.801 0.569 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.380 0.348 0.492 0.543 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.800 0.693 4.011 0.776 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.355 0.296 4.356 0.761 ;
      RECT 4.339 0.296 4.355 0.973 ;
      RECT 4.295 0.296 4.339 1.021 ;
      RECT 4.056 0.296 4.295 0.351 ;
      RECT 4.281 0.706 4.295 1.021 ;
      RECT 4.248 0.829 4.281 1.021 ;
      RECT 3.995 0.174 4.056 0.351 ;
      RECT 3.965 0.174 3.995 0.255 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.035 0.417 1.195 0.502 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.168 0.517 0.295 0.627 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.248 -0.080 4.400 0.080 ;
      RECT 4.157 -0.080 4.248 0.211 ;
      RECT 3.852 -0.080 4.157 0.080 ;
      RECT 3.601 -0.080 3.852 0.122 ;
      RECT 3.297 -0.080 3.601 0.080 ;
      RECT 3.207 -0.080 3.297 0.122 ;
      RECT 2.516 -0.080 3.207 0.080 ;
      RECT 2.425 -0.080 2.516 0.254 ;
      RECT 1.776 -0.080 2.425 0.080 ;
      RECT 1.685 -0.080 1.776 0.327 ;
      RECT 0.837 -0.080 1.685 0.080 ;
      RECT 0.747 -0.080 0.837 0.122 ;
      RECT 0.288 -0.080 0.747 0.080 ;
      RECT 0.197 -0.080 0.288 0.122 ;
      RECT 0.000 -0.080 0.197 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.997 1.120 4.400 1.280 ;
      RECT 3.907 0.857 3.997 1.280 ;
      RECT 3.395 1.120 3.907 1.280 ;
      RECT 3.284 1.078 3.395 1.280 ;
      RECT 2.628 1.120 3.284 1.280 ;
      RECT 2.517 1.078 2.628 1.280 ;
      RECT 1.781 1.120 2.517 1.280 ;
      RECT 1.691 0.963 1.781 1.280 ;
      RECT 0.933 1.120 1.691 1.280 ;
      RECT 0.843 1.001 0.933 1.280 ;
      RECT 0.245 1.120 0.843 1.280 ;
      RECT 0.155 0.932 0.245 1.280 ;
      RECT 0.000 1.120 0.155 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.093 0.407 4.184 0.488 ;
      RECT 3.840 0.407 4.093 0.462 ;
      RECT 3.679 0.583 4.088 0.638 ;
      RECT 3.779 0.206 3.840 0.462 ;
      RECT 3.713 0.952 3.804 1.033 ;
      RECT 3.393 0.206 3.779 0.261 ;
      RECT 3.559 0.952 3.713 1.020 ;
      RECT 3.679 0.327 3.692 0.408 ;
      RECT 3.617 0.327 3.679 0.638 ;
      RECT 3.601 0.327 3.617 0.408 ;
      RECT 3.559 0.526 3.617 0.638 ;
      RECT 3.527 0.526 3.559 1.020 ;
      RECT 3.497 0.573 3.527 1.020 ;
      RECT 2.247 0.939 3.497 0.994 ;
      RECT 3.388 0.336 3.479 0.417 ;
      RECT 3.295 0.206 3.393 0.273 ;
      RECT 3.360 0.362 3.388 0.417 ;
      RECT 3.299 0.362 3.360 0.833 ;
      RECT 3.269 0.614 3.299 0.833 ;
      RECT 3.141 0.206 3.295 0.261 ;
      RECT 3.211 0.614 3.269 0.695 ;
      RECT 3.080 0.206 3.141 0.857 ;
      RECT 2.933 0.206 3.080 0.263 ;
      RECT 3.016 0.802 3.080 0.857 ;
      RECT 2.965 0.382 3.017 0.463 ;
      RECT 2.925 0.802 3.016 0.883 ;
      RECT 2.927 0.382 2.965 0.727 ;
      RECT 2.857 0.206 2.933 0.304 ;
      RECT 2.904 0.395 2.927 0.727 ;
      RECT 2.843 0.223 2.857 0.304 ;
      RECT 2.781 0.380 2.843 0.883 ;
      RECT 2.780 0.380 2.781 0.435 ;
      RECT 2.733 0.802 2.781 0.883 ;
      RECT 2.720 0.267 2.780 0.435 ;
      RECT 2.719 0.240 2.720 0.435 ;
      RECT 2.657 0.548 2.720 0.644 ;
      RECT 2.629 0.240 2.719 0.321 ;
      RECT 2.596 0.390 2.657 0.852 ;
      RECT 2.384 0.390 2.596 0.445 ;
      RECT 2.472 0.798 2.596 0.852 ;
      RECT 2.473 0.501 2.535 0.694 ;
      RECT 1.987 0.501 2.473 0.556 ;
      RECT 2.381 0.798 2.472 0.879 ;
      RECT 2.348 0.364 2.384 0.445 ;
      RECT 2.287 0.163 2.348 0.445 ;
      RECT 1.856 0.163 2.287 0.218 ;
      RECT 2.213 0.627 2.247 0.994 ;
      RECT 2.185 0.614 2.213 0.994 ;
      RECT 2.123 0.614 2.185 0.695 ;
      RECT 1.949 0.411 1.987 0.876 ;
      RECT 1.925 0.398 1.949 0.876 ;
      RECT 1.859 0.398 1.925 0.479 ;
      RECT 1.880 0.795 1.925 0.876 ;
      RECT 1.803 0.614 1.864 0.701 ;
      RECT 1.672 0.424 1.859 0.479 ;
      RECT 1.476 0.646 1.803 0.701 ;
      RECT 1.611 0.424 1.672 0.564 ;
      RECT 1.581 0.483 1.611 0.564 ;
      RECT 1.459 0.890 1.549 0.971 ;
      RECT 1.449 0.249 1.476 0.701 ;
      RECT 1.319 0.890 1.459 0.945 ;
      RECT 1.415 0.249 1.449 0.792 ;
      RECT 1.413 0.249 1.415 0.304 ;
      RECT 1.388 0.646 1.415 0.792 ;
      RECT 1.323 0.223 1.413 0.304 ;
      RECT 1.257 0.436 1.319 0.945 ;
      RECT 0.613 0.732 1.257 0.787 ;
      RECT 1.109 0.206 1.200 0.293 ;
      RECT 1.135 0.856 1.196 0.962 ;
      RECT 0.736 0.856 1.135 0.911 ;
      RECT 0.475 0.206 1.109 0.261 ;
      RECT 0.911 0.317 0.912 0.398 ;
      RECT 0.821 0.317 0.911 0.402 ;
      RECT 0.649 0.348 0.821 0.402 ;
      RECT 0.675 0.856 0.736 0.993 ;
      RECT 0.649 0.595 0.691 0.676 ;
      RECT 0.624 0.938 0.675 0.993 ;
      RECT 0.600 0.348 0.649 0.676 ;
      RECT 0.533 0.938 0.624 1.019 ;
      RECT 0.552 0.732 0.613 0.860 ;
      RECT 0.572 0.348 0.600 0.663 ;
      RECT 0.557 0.348 0.572 0.429 ;
      RECT 0.491 0.608 0.572 0.663 ;
      RECT 0.139 0.805 0.552 0.860 ;
      RECT 0.429 0.608 0.491 0.748 ;
      RECT 0.384 0.152 0.475 0.261 ;
      RECT 0.400 0.667 0.429 0.748 ;
      RECT 0.105 0.317 0.139 0.398 ;
      RECT 0.105 0.688 0.139 0.860 ;
      RECT 0.077 0.317 0.105 0.860 ;
      RECT 0.044 0.317 0.077 0.769 ;
  END
END SDFFRHQX1

MACRO SDFFRXL
  CLASS CORE ;
  FOREIGN SDFFRXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.974 0.552 1.005 0.637 ;
      RECT 0.884 0.552 0.974 0.696 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.325 0.429 0.480 0.545 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.928 0.690 2.018 0.771 ;
      RECT 1.888 0.690 1.928 0.767 ;
      RECT 1.868 0.562 1.888 0.767 ;
      RECT 1.827 0.562 1.868 0.758 ;
      RECT 1.792 0.562 1.827 0.638 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.445 0.206 4.506 0.961 ;
      RECT 4.351 0.206 4.445 0.261 ;
      RECT 4.405 0.833 4.445 0.961 ;
      RECT 4.372 0.906 4.405 0.961 ;
      RECT 4.282 0.906 4.372 1.007 ;
      RECT 4.261 0.151 4.351 0.261 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.809 0.862 4.831 0.943 ;
      RECT 4.748 0.450 4.809 0.943 ;
      RECT 4.725 0.450 4.748 0.505 ;
      RECT 4.741 0.862 4.748 0.943 ;
      RECT 4.587 0.283 4.725 0.505 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.088 0.375 1.192 0.501 ;
      RECT 1.070 0.408 1.088 0.495 ;
      RECT 1.055 0.414 1.070 0.495 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.167 0.646 0.313 0.767 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.545 -0.080 4.900 0.080 ;
      RECT 4.455 -0.080 4.545 0.122 ;
      RECT 4.118 -0.080 4.455 0.080 ;
      RECT 4.028 -0.080 4.118 0.211 ;
      RECT 3.651 -0.080 4.028 0.080 ;
      RECT 3.561 -0.080 3.651 0.249 ;
      RECT 2.388 -0.080 3.561 0.080 ;
      RECT 2.793 0.302 2.884 0.404 ;
      RECT 2.466 0.302 2.793 0.352 ;
      RECT 2.388 0.302 2.466 0.361 ;
      RECT 2.327 -0.080 2.388 0.361 ;
      RECT 1.853 -0.080 2.327 0.080 ;
      RECT 1.763 -0.080 1.853 0.214 ;
      RECT 0.875 -0.080 1.763 0.080 ;
      RECT 0.785 -0.080 0.875 0.122 ;
      RECT 0.321 -0.080 0.785 0.080 ;
      RECT 0.231 -0.080 0.321 0.122 ;
      RECT 0.000 -0.080 0.231 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.627 1.120 4.900 1.280 ;
      RECT 4.537 1.078 4.627 1.280 ;
      RECT 4.171 1.120 4.537 1.280 ;
      RECT 4.081 0.989 4.171 1.280 ;
      RECT 3.634 1.120 4.081 1.280 ;
      RECT 3.544 0.986 3.634 1.280 ;
      RECT 3.015 1.120 3.544 1.280 ;
      RECT 2.766 0.986 3.015 1.280 ;
      RECT 1.954 1.120 2.766 1.280 ;
      RECT 1.864 1.078 1.954 1.280 ;
      RECT 0.989 1.120 1.864 1.280 ;
      RECT 0.899 0.986 0.989 1.280 ;
      RECT 0.202 1.120 0.899 1.280 ;
      RECT 0.111 1.078 0.202 1.280 ;
      RECT 0.000 1.120 0.111 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.343 0.329 4.372 0.752 ;
      RECT 4.282 0.329 4.343 0.798 ;
      RECT 4.234 0.329 4.282 0.440 ;
      RECT 4.253 0.671 4.282 0.798 ;
      RECT 4.143 0.448 4.155 0.529 ;
      RECT 4.140 0.444 4.143 0.529 ;
      RECT 4.008 0.444 4.140 0.535 ;
      RECT 3.947 0.444 4.008 0.917 ;
      RECT 3.891 0.444 3.947 0.499 ;
      RECT 3.821 0.862 3.947 0.917 ;
      RECT 3.830 0.218 3.891 0.499 ;
      RECT 3.794 0.715 3.884 0.807 ;
      RECT 3.788 0.218 3.830 0.435 ;
      RECT 3.731 0.862 3.821 0.943 ;
      RECT 3.493 0.752 3.794 0.807 ;
      RECT 3.694 0.380 3.788 0.435 ;
      RECT 3.633 0.380 3.694 0.614 ;
      RECT 3.603 0.533 3.633 0.614 ;
      RECT 3.446 0.333 3.493 0.811 ;
      RECT 3.446 0.952 3.447 1.033 ;
      RECT 3.432 0.333 3.446 1.033 ;
      RECT 3.243 0.333 3.432 0.388 ;
      RECT 3.385 0.752 3.432 1.033 ;
      RECT 3.357 0.952 3.385 1.033 ;
      RECT 3.325 0.569 3.340 0.650 ;
      RECT 3.249 0.569 3.325 0.685 ;
      RECT 3.228 0.630 3.249 0.685 ;
      RECT 3.153 0.307 3.243 0.388 ;
      RECT 3.167 0.630 3.228 0.917 ;
      RECT 2.783 0.862 3.167 0.917 ;
      RECT 3.069 0.485 3.150 0.565 ;
      RECT 3.008 0.161 3.069 0.806 ;
      RECT 2.564 0.161 3.008 0.215 ;
      RECT 2.845 0.751 3.008 0.806 ;
      RECT 2.549 0.510 2.925 0.590 ;
      RECT 2.722 0.669 2.783 0.917 ;
      RECT 2.687 0.862 2.722 0.917 ;
      RECT 2.626 0.862 2.687 1.039 ;
      RECT 2.076 0.985 2.626 1.039 ;
      RECT 2.474 0.151 2.564 0.232 ;
      RECT 2.488 0.435 2.549 0.879 ;
      RECT 2.237 0.435 2.488 0.489 ;
      RECT 2.408 0.824 2.488 0.879 ;
      RECT 2.317 0.824 2.408 0.905 ;
      RECT 2.315 0.581 2.405 0.662 ;
      RECT 2.198 0.594 2.315 0.649 ;
      RECT 2.176 0.262 2.237 0.489 ;
      RECT 2.137 0.580 2.198 0.921 ;
      RECT 2.146 0.262 2.176 0.449 ;
      RECT 1.734 0.394 2.146 0.449 ;
      RECT 2.093 0.580 2.137 0.635 ;
      RECT 2.003 0.504 2.093 0.635 ;
      RECT 2.015 0.954 2.076 1.039 ;
      RECT 1.998 0.183 2.070 0.264 ;
      RECT 1.762 0.954 2.015 1.008 ;
      RECT 1.979 0.183 1.998 0.338 ;
      RECT 1.937 0.196 1.979 0.338 ;
      RECT 1.574 0.283 1.937 0.338 ;
      RECT 1.722 0.954 1.762 1.037 ;
      RECT 1.644 0.394 1.734 0.495 ;
      RECT 1.701 0.954 1.722 1.050 ;
      RECT 1.632 0.969 1.701 1.050 ;
      RECT 1.491 0.982 1.632 1.037 ;
      RECT 1.574 0.596 1.613 0.905 ;
      RECT 1.552 0.283 1.574 0.905 ;
      RECT 1.513 0.283 1.552 0.651 ;
      RECT 1.458 0.283 1.513 0.338 ;
      RECT 1.430 0.707 1.491 1.037 ;
      RECT 1.368 0.233 1.458 0.338 ;
      RECT 1.379 0.707 1.430 0.762 ;
      RECT 1.134 0.982 1.430 1.037 ;
      RECT 1.350 0.463 1.379 0.762 ;
      RECT 1.309 0.824 1.370 0.905 ;
      RECT 1.318 0.450 1.350 0.762 ;
      RECT 1.259 0.450 1.318 0.531 ;
      RECT 1.257 0.824 1.309 0.879 ;
      RECT 1.196 0.752 1.257 0.879 ;
      RECT 1.212 0.229 1.236 0.310 ;
      RECT 1.145 0.206 1.212 0.310 ;
      RECT 0.719 0.752 1.196 0.807 ;
      RECT 0.571 0.206 1.145 0.261 ;
      RECT 1.073 0.862 1.134 1.037 ;
      RECT 0.837 0.862 1.073 0.917 ;
      RECT 0.841 0.385 0.931 0.465 ;
      RECT 0.644 0.398 0.841 0.452 ;
      RECT 0.776 0.862 0.837 1.006 ;
      RECT 0.370 0.951 0.776 1.006 ;
      RECT 0.628 0.726 0.719 0.807 ;
      RECT 0.630 0.345 0.644 0.452 ;
      RECT 0.630 0.590 0.631 0.671 ;
      RECT 0.569 0.345 0.630 0.671 ;
      RECT 0.514 0.163 0.571 0.261 ;
      RECT 0.554 0.345 0.569 0.426 ;
      RECT 0.541 0.590 0.569 0.671 ;
      RECT 0.513 0.617 0.541 0.671 ;
      RECT 0.513 0.815 0.528 0.896 ;
      RECT 0.510 0.150 0.514 0.261 ;
      RECT 0.452 0.617 0.513 0.896 ;
      RECT 0.424 0.150 0.510 0.231 ;
      RECT 0.437 0.815 0.452 0.896 ;
      RECT 0.309 0.892 0.370 1.006 ;
      RECT 0.143 0.892 0.309 0.946 ;
      RECT 0.105 0.293 0.143 0.374 ;
      RECT 0.105 0.840 0.143 0.946 ;
      RECT 0.044 0.293 0.105 0.946 ;
  END
END SDFFRXL

MACRO SDFFRX4
  CLASS CORE ;
  FOREIGN SDFFRX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.746 0.488 0.836 0.663 ;
      RECT 0.734 0.490 0.746 0.663 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.466 0.307 0.470 0.557 ;
      RECT 0.388 0.306 0.466 0.557 ;
      RECT 0.378 0.306 0.388 0.548 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.933 0.654 2.054 0.832 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.440 0.285 5.540 0.767 ;
      RECT 5.435 0.285 5.440 0.365 ;
      RECT 5.435 0.662 5.440 0.743 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.862 0.300 5.889 0.743 ;
      RECT 5.788 0.285 5.862 0.743 ;
      RECT 5.787 0.285 5.788 0.494 ;
      RECT 5.773 0.662 5.788 0.743 ;
      RECT 5.773 0.285 5.787 0.365 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.042 0.562 1.102 0.643 ;
      RECT 1.007 0.562 1.042 0.617 ;
      RECT 0.947 0.439 1.007 0.617 ;
      RECT 0.928 0.439 0.947 0.494 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.174 0.560 0.296 0.675 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.031 -0.080 6.100 0.080 ;
      RECT 5.942 -0.080 6.031 0.211 ;
      RECT 5.693 -0.080 5.942 0.080 ;
      RECT 5.604 -0.080 5.693 0.211 ;
      RECT 5.355 -0.080 5.604 0.080 ;
      RECT 5.266 -0.080 5.355 0.211 ;
      RECT 4.994 -0.080 5.266 0.080 ;
      RECT 4.904 -0.080 4.994 0.211 ;
      RECT 4.613 -0.080 4.904 0.080 ;
      RECT 4.524 -0.080 4.613 0.211 ;
      RECT 4.228 -0.080 4.524 0.080 ;
      RECT 4.138 -0.080 4.228 0.211 ;
      RECT 3.760 -0.080 4.138 0.080 ;
      RECT 3.671 -0.080 3.760 0.242 ;
      RECT 3.075 -0.080 3.671 0.080 ;
      RECT 3.014 -0.080 3.075 0.336 ;
      RECT 2.585 -0.080 3.014 0.080 ;
      RECT 2.495 -0.080 2.585 0.214 ;
      RECT 2.054 -0.080 2.495 0.080 ;
      RECT 1.965 -0.080 2.054 0.303 ;
      RECT 0.856 -0.080 1.965 0.080 ;
      RECT 0.766 -0.080 0.856 0.122 ;
      RECT 0.285 -0.080 0.766 0.080 ;
      RECT 0.195 -0.080 0.285 0.122 ;
      RECT 0.000 -0.080 0.195 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.031 1.120 6.100 1.280 ;
      RECT 5.942 0.977 6.031 1.280 ;
      RECT 5.693 1.120 5.942 1.280 ;
      RECT 5.604 0.977 5.693 1.280 ;
      RECT 5.355 1.120 5.604 1.280 ;
      RECT 5.266 0.986 5.355 1.280 ;
      RECT 4.941 1.120 5.266 1.280 ;
      RECT 4.851 0.742 4.941 1.280 ;
      RECT 4.254 1.120 4.851 1.280 ;
      RECT 4.164 0.986 4.254 1.280 ;
      RECT 3.599 1.120 4.164 1.280 ;
      RECT 3.509 0.890 3.599 1.280 ;
      RECT 2.847 1.120 3.509 1.280 ;
      RECT 2.757 0.948 2.847 1.280 ;
      RECT 1.880 1.120 2.757 1.280 ;
      RECT 1.790 1.078 1.880 1.280 ;
      RECT 1.025 1.120 1.790 1.280 ;
      RECT 0.935 0.986 1.025 1.280 ;
      RECT 0.224 1.120 0.935 1.280 ;
      RECT 0.135 1.078 0.224 1.280 ;
      RECT 0.000 1.120 0.135 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.969 0.483 6.030 0.893 ;
      RECT 5.354 0.838 5.969 0.893 ;
      RECT 5.293 0.332 5.354 0.893 ;
      RECT 5.173 0.332 5.293 0.412 ;
      RECT 5.131 0.777 5.293 0.832 ;
      RECT 4.967 0.500 5.215 0.581 ;
      RECT 5.083 0.331 5.173 0.412 ;
      RECT 5.041 0.708 5.131 0.901 ;
      RECT 5.081 0.332 5.083 0.399 ;
      RECT 4.803 0.513 4.967 0.568 ;
      RECT 4.743 0.171 4.803 0.640 ;
      RECT 4.714 0.171 4.743 0.351 ;
      RECT 4.603 0.586 4.743 0.640 ;
      RECT 4.423 0.296 4.714 0.351 ;
      RECT 4.583 0.411 4.677 0.492 ;
      RECT 4.542 0.586 4.603 0.913 ;
      RECT 4.428 0.411 4.583 0.501 ;
      RECT 4.513 0.711 4.542 0.913 ;
      RECT 4.093 0.858 4.513 0.913 ;
      RECT 4.163 0.446 4.428 0.501 ;
      RECT 4.362 0.167 4.423 0.351 ;
      RECT 4.333 0.167 4.362 0.248 ;
      RECT 4.102 0.356 4.163 0.801 ;
      RECT 3.484 0.356 4.102 0.413 ;
      RECT 3.936 0.746 4.102 0.801 ;
      RECT 4.032 0.858 4.093 1.012 ;
      RECT 3.899 0.577 3.989 0.671 ;
      RECT 3.936 0.893 3.950 0.974 ;
      RECT 3.875 0.746 3.936 0.974 ;
      RECT 3.363 0.577 3.899 0.632 ;
      RECT 3.432 0.746 3.875 0.801 ;
      RECT 3.861 0.893 3.875 0.974 ;
      RECT 3.424 0.261 3.484 0.413 ;
      RECT 3.371 0.746 3.432 0.918 ;
      RECT 3.314 0.261 3.424 0.315 ;
      RECT 3.261 0.863 3.371 0.918 ;
      RECT 3.302 0.414 3.363 0.632 ;
      RECT 3.227 0.577 3.302 0.632 ;
      RECT 3.171 0.863 3.261 0.950 ;
      RECT 3.166 0.415 3.227 0.749 ;
      RECT 2.843 0.415 3.166 0.470 ;
      RECT 3.049 0.694 3.166 0.749 ;
      RECT 2.687 0.531 3.105 0.586 ;
      RECT 3.047 0.694 3.049 0.939 ;
      RECT 2.988 0.694 3.047 0.952 ;
      RECT 2.958 0.871 2.988 0.952 ;
      RECT 2.853 0.676 2.897 0.757 ;
      RECT 2.793 0.676 2.853 0.871 ;
      RECT 2.782 0.161 2.843 0.470 ;
      RECT 2.653 0.817 2.793 0.871 ;
      RECT 2.651 0.161 2.782 0.215 ;
      RECT 2.626 0.373 2.687 0.749 ;
      RECT 2.592 0.817 2.653 1.039 ;
      RECT 2.437 0.373 2.626 0.427 ;
      RECT 2.509 0.694 2.626 0.749 ;
      RECT 2.024 0.985 2.592 1.039 ;
      RECT 2.419 0.694 2.509 0.921 ;
      RECT 2.411 0.500 2.501 0.581 ;
      RECT 2.348 0.340 2.437 0.427 ;
      RECT 2.196 0.513 2.411 0.568 ;
      RECT 1.838 0.373 2.348 0.427 ;
      RECT 2.196 0.848 2.210 0.929 ;
      RECT 2.135 0.482 2.196 0.929 ;
      RECT 1.999 0.482 2.135 0.537 ;
      RECT 2.120 0.848 2.135 0.929 ;
      RECT 1.963 0.939 2.024 1.039 ;
      RECT 1.707 0.939 1.963 0.994 ;
      RECT 1.777 0.373 1.838 0.633 ;
      RECT 1.485 0.196 1.835 0.251 ;
      RECT 1.748 0.552 1.777 0.633 ;
      RECT 1.666 0.723 1.707 1.035 ;
      RECT 1.646 0.471 1.666 1.035 ;
      RECT 1.606 0.471 1.646 0.777 ;
      RECT 1.153 0.980 1.646 1.035 ;
      RECT 1.345 0.471 1.606 0.526 ;
      RECT 1.496 0.833 1.563 0.914 ;
      RECT 1.435 0.587 1.496 0.914 ;
      RECT 1.426 0.196 1.485 0.337 ;
      RECT 1.224 0.587 1.435 0.642 ;
      RECT 1.425 0.196 1.426 0.350 ;
      RECT 1.411 0.269 1.425 0.350 ;
      RECT 1.336 0.269 1.411 0.389 ;
      RECT 1.327 0.817 1.373 0.898 ;
      RECT 1.285 0.445 1.345 0.526 ;
      RECT 1.224 0.335 1.336 0.389 ;
      RECT 1.266 0.746 1.327 0.898 ;
      RECT 0.729 0.746 1.266 0.801 ;
      RECT 1.163 0.335 1.224 0.642 ;
      RECT 1.125 0.198 1.215 0.279 ;
      RECT 1.092 0.861 1.153 1.035 ;
      RECT 0.691 0.206 1.125 0.261 ;
      RECT 0.856 0.861 1.092 0.915 ;
      RECT 0.654 0.320 0.930 0.375 ;
      RECT 0.795 0.861 0.856 1.008 ;
      RECT 0.137 0.954 0.795 1.008 ;
      RECT 0.654 0.746 0.729 0.857 ;
      RECT 0.630 0.162 0.691 0.261 ;
      RECT 0.566 0.320 0.654 0.677 ;
      RECT 0.639 0.776 0.654 0.857 ;
      RECT 0.407 0.162 0.630 0.217 ;
      RECT 0.547 0.324 0.566 0.405 ;
      RECT 0.556 0.623 0.566 0.677 ;
      RECT 0.495 0.623 0.556 0.869 ;
      RECT 0.486 0.814 0.495 0.869 ;
      RECT 0.396 0.814 0.486 0.895 ;
      RECT 0.107 0.301 0.137 0.382 ;
      RECT 0.107 0.757 0.137 1.008 ;
      RECT 0.077 0.301 0.107 1.008 ;
      RECT 0.046 0.301 0.077 0.838 ;
  END
END SDFFRX4

MACRO SDFFNRX1
  CLASS CORE ;
  FOREIGN SDFFNRX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.886 0.560 1.008 0.681 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.324 0.419 0.477 0.529 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.890 0.795 2.056 0.850 ;
      RECT 1.829 0.569 1.890 0.850 ;
      RECT 1.786 0.569 1.829 0.631 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.489 0.205 4.497 0.785 ;
      RECT 4.436 0.205 4.489 0.900 ;
      RECT 4.389 0.205 4.436 0.306 ;
      RECT 4.409 0.730 4.436 0.900 ;
      RECT 4.320 0.839 4.409 0.900 ;
      RECT 4.204 0.205 4.389 0.260 ;
      RECT 4.260 0.839 4.320 0.950 ;
      RECT 4.220 0.869 4.260 0.950 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.653 0.302 4.656 0.871 ;
      RECT 4.588 0.302 4.653 0.937 ;
      RECT 4.583 0.302 4.588 0.439 ;
      RECT 4.563 0.744 4.588 0.937 ;
      RECT 4.563 0.323 4.583 0.439 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.060 0.381 1.166 0.505 ;
      RECT 1.039 0.385 1.060 0.505 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.166 0.636 0.311 0.769 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.631 -0.080 4.700 0.080 ;
      RECT 4.542 -0.080 4.631 0.122 ;
      RECT 3.927 -0.080 4.542 0.080 ;
      RECT 3.838 -0.080 3.927 0.122 ;
      RECT 3.526 -0.080 3.838 0.080 ;
      RECT 3.437 -0.080 3.526 0.122 ;
      RECT 2.375 -0.080 3.437 0.080 ;
      RECT 2.843 0.358 2.872 0.409 ;
      RECT 2.783 0.302 2.843 0.409 ;
      RECT 2.453 0.302 2.783 0.352 ;
      RECT 2.375 0.302 2.453 0.352 ;
      RECT 2.314 -0.080 2.375 0.352 ;
      RECT 1.844 -0.080 2.314 0.080 ;
      RECT 1.754 -0.080 1.844 0.214 ;
      RECT 0.844 -0.080 1.754 0.080 ;
      RECT 0.754 -0.080 0.844 0.122 ;
      RECT 0.142 -0.080 0.754 0.080 ;
      RECT 0.053 -0.080 0.142 0.122 ;
      RECT 0.000 -0.080 0.053 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.629 1.120 4.700 1.280 ;
      RECT 4.513 1.078 4.629 1.280 ;
      RECT 4.120 1.120 4.513 1.280 ;
      RECT 4.030 0.877 4.120 1.280 ;
      RECT 3.598 1.120 4.030 1.280 ;
      RECT 3.508 0.984 3.598 1.280 ;
      RECT 2.999 1.120 3.508 1.280 ;
      RECT 2.751 0.984 2.999 1.280 ;
      RECT 1.925 1.120 2.751 1.280 ;
      RECT 1.836 1.078 1.925 1.280 ;
      RECT 0.984 1.120 1.836 1.280 ;
      RECT 0.894 0.986 0.984 1.280 ;
      RECT 0.298 1.120 0.894 1.280 ;
      RECT 0.208 1.078 0.298 1.280 ;
      RECT 0.000 1.120 0.208 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.316 0.512 4.331 0.593 ;
      RECT 4.281 0.511 4.316 0.593 ;
      RECT 4.203 0.511 4.281 0.740 ;
      RECT 4.191 0.314 4.203 0.740 ;
      RECT 4.142 0.314 4.191 0.565 ;
      RECT 4.072 0.314 4.142 0.369 ;
      RECT 4.021 0.435 4.082 0.785 ;
      RECT 3.983 0.288 4.072 0.369 ;
      RECT 3.906 0.435 4.021 0.489 ;
      RECT 3.782 0.730 4.021 0.785 ;
      RECT 3.845 0.380 3.906 0.489 ;
      RECT 3.727 0.380 3.845 0.435 ;
      RECT 3.695 0.510 3.785 0.590 ;
      RECT 3.721 0.730 3.782 0.908 ;
      RECT 3.637 0.162 3.727 0.435 ;
      RECT 3.692 0.827 3.721 0.908 ;
      RECT 3.384 0.535 3.695 0.589 ;
      RECT 3.547 0.380 3.637 0.435 ;
      RECT 3.458 0.380 3.547 0.480 ;
      RECT 3.384 0.952 3.413 1.033 ;
      RECT 3.323 0.481 3.384 1.033 ;
      RECT 3.206 0.481 3.323 0.536 ;
      RECT 3.215 0.158 3.305 0.239 ;
      RECT 3.197 0.595 3.226 0.676 ;
      RECT 3.206 0.312 3.220 0.393 ;
      RECT 3.053 0.161 3.215 0.215 ;
      RECT 3.145 0.312 3.206 0.536 ;
      RECT 3.136 0.595 3.197 0.793 ;
      RECT 3.131 0.312 3.145 0.393 ;
      RECT 3.053 0.738 3.136 0.793 ;
      RECT 2.992 0.161 3.053 0.793 ;
      RECT 2.525 0.161 2.992 0.215 ;
      RECT 2.889 0.738 2.992 0.793 ;
      RECT 2.819 0.481 2.909 0.574 ;
      RECT 2.829 0.738 2.889 0.851 ;
      RECT 2.536 0.519 2.819 0.574 ;
      RECT 2.707 0.644 2.768 0.911 ;
      RECT 2.673 0.856 2.707 0.911 ;
      RECT 2.612 0.856 2.673 1.039 ;
      RECT 2.047 0.985 2.612 1.039 ;
      RECT 2.475 0.435 2.536 0.806 ;
      RECT 2.436 0.151 2.525 0.232 ;
      RECT 2.238 0.435 2.475 0.489 ;
      RECT 2.395 0.751 2.475 0.806 ;
      RECT 2.334 0.751 2.395 0.910 ;
      RECT 2.303 0.581 2.392 0.662 ;
      RECT 2.305 0.829 2.334 0.910 ;
      RECT 2.196 0.594 2.303 0.649 ;
      RECT 2.177 0.265 2.238 0.489 ;
      RECT 2.196 0.829 2.210 0.910 ;
      RECT 2.135 0.580 2.196 0.910 ;
      RECT 2.130 0.265 2.177 0.449 ;
      RECT 2.081 0.580 2.135 0.635 ;
      RECT 2.121 0.829 2.135 0.910 ;
      RECT 1.725 0.394 2.130 0.449 ;
      RECT 1.985 0.505 2.081 0.635 ;
      RECT 1.987 0.183 2.065 0.264 ;
      RECT 1.986 0.939 2.047 1.039 ;
      RECT 1.927 0.183 1.987 0.338 ;
      RECT 1.753 0.939 1.986 0.994 ;
      RECT 1.451 0.283 1.927 0.338 ;
      RECT 1.697 0.699 1.753 1.029 ;
      RECT 1.635 0.394 1.725 0.495 ;
      RECT 1.692 0.570 1.697 1.029 ;
      RECT 1.637 0.570 1.692 0.754 ;
      RECT 1.128 0.974 1.692 1.029 ;
      RECT 1.550 0.570 1.637 0.625 ;
      RECT 1.515 0.829 1.604 0.914 ;
      RECT 1.489 0.462 1.550 0.625 ;
      RECT 1.455 0.680 1.515 0.914 ;
      RECT 1.445 0.462 1.489 0.543 ;
      RECT 1.408 0.680 1.455 0.735 ;
      RECT 1.362 0.276 1.451 0.357 ;
      RECT 1.362 0.617 1.408 0.735 ;
      RECT 1.295 0.818 1.385 0.905 ;
      RECT 1.348 0.276 1.362 0.735 ;
      RECT 1.302 0.276 1.348 0.671 ;
      RECT 1.265 0.818 1.295 0.873 ;
      RECT 1.204 0.738 1.265 0.873 ;
      RECT 0.720 0.738 1.204 0.793 ;
      RECT 1.113 0.206 1.203 0.298 ;
      RECT 1.067 0.862 1.128 1.029 ;
      RECT 0.568 0.206 1.113 0.261 ;
      RECT 0.823 0.862 1.067 0.917 ;
      RECT 0.836 0.317 0.926 0.398 ;
      RECT 0.641 0.330 0.836 0.385 ;
      RECT 0.762 0.862 0.823 0.946 ;
      RECT 0.145 0.892 0.762 0.946 ;
      RECT 0.630 0.725 0.720 0.806 ;
      RECT 0.626 0.586 0.680 0.667 ;
      RECT 0.626 0.330 0.641 0.417 ;
      RECT 0.591 0.330 0.626 0.667 ;
      RECT 0.566 0.330 0.591 0.654 ;
      RECT 0.508 0.158 0.568 0.261 ;
      RECT 0.551 0.330 0.566 0.417 ;
      RECT 0.525 0.599 0.566 0.654 ;
      RECT 0.464 0.599 0.525 0.771 ;
      RECT 0.396 0.158 0.508 0.213 ;
      RECT 0.435 0.690 0.464 0.771 ;
      RECT 0.104 0.838 0.145 0.946 ;
      RECT 0.104 0.321 0.142 0.402 ;
      RECT 0.044 0.321 0.104 0.946 ;
  END
END SDFFNRX1

MACRO SDFFNXL
  CLASS CORE ;
  FOREIGN SDFFNXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.719 0.433 0.844 0.500 ;
      RECT 0.631 0.412 0.719 0.500 ;
      RECT 0.617 0.412 0.631 0.467 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.978 0.619 1.069 0.700 ;
      RECT 0.849 0.632 0.978 0.687 ;
      RECT 0.788 0.567 0.849 0.687 ;
      RECT 0.566 0.567 0.788 0.633 ;
      RECT 0.531 0.573 0.566 0.627 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.470 0.837 3.561 0.918 ;
      RECT 3.466 0.292 3.476 0.373 ;
      RECT 3.466 0.837 3.470 0.894 ;
      RECT 3.405 0.292 3.466 0.892 ;
      RECT 3.385 0.292 3.405 0.373 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.137 0.150 3.227 0.249 ;
      RECT 3.127 0.487 3.178 0.819 ;
      RECT 3.110 0.194 3.137 0.249 ;
      RECT 3.117 0.487 3.127 0.845 ;
      RECT 3.110 0.487 3.117 0.542 ;
      RECT 3.037 0.764 3.117 0.845 ;
      RECT 3.049 0.194 3.110 0.542 ;
      RECT 2.876 0.306 3.049 0.361 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.133 0.439 1.176 0.494 ;
      RECT 1.057 0.335 1.133 0.494 ;
      RECT 1.042 0.335 1.057 0.415 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.234 0.537 0.315 0.633 ;
      RECT 0.214 0.524 0.234 0.633 ;
      RECT 0.172 0.524 0.214 0.632 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.448 -0.080 3.700 0.080 ;
      RECT 3.357 -0.080 3.448 0.122 ;
      RECT 3.025 -0.080 3.357 0.080 ;
      RECT 2.934 -0.080 3.025 0.122 ;
      RECT 2.373 -0.080 2.934 0.080 ;
      RECT 2.282 -0.080 2.373 0.345 ;
      RECT 1.745 -0.080 2.282 0.080 ;
      RECT 1.683 -0.080 1.745 0.259 ;
      RECT 0.820 -0.080 1.683 0.080 ;
      RECT 0.729 -0.080 0.820 0.122 ;
      RECT 0.304 -0.080 0.729 0.080 ;
      RECT 0.304 0.322 0.352 0.373 ;
      RECT 0.262 -0.080 0.304 0.373 ;
      RECT 0.243 -0.080 0.262 0.360 ;
      RECT 0.000 -0.080 0.243 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.341 1.120 3.700 1.280 ;
      RECT 3.250 1.065 3.341 1.280 ;
      RECT 2.914 1.120 3.250 1.280 ;
      RECT 2.823 1.078 2.914 1.280 ;
      RECT 2.193 1.120 2.823 1.280 ;
      RECT 1.851 1.078 2.193 1.280 ;
      RECT 1.069 1.120 1.851 1.280 ;
      RECT 0.978 1.065 1.069 1.280 ;
      RECT 0.251 1.120 0.978 1.280 ;
      RECT 0.141 1.078 0.251 1.280 ;
      RECT 0.000 1.120 0.141 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.262 0.337 3.324 0.995 ;
      RECT 3.171 0.324 3.262 0.405 ;
      RECT 3.133 0.940 3.262 0.995 ;
      RECT 3.071 0.940 3.133 1.036 ;
      RECT 3.013 0.954 3.071 1.036 ;
      RECT 2.985 0.623 3.053 0.704 ;
      RECT 2.815 0.954 3.013 1.008 ;
      RECT 2.962 0.538 2.985 0.704 ;
      RECT 2.923 0.538 2.962 0.677 ;
      RECT 2.715 0.538 2.923 0.593 ;
      RECT 2.513 0.189 2.822 0.244 ;
      RECT 2.754 0.654 2.815 1.008 ;
      RECT 2.724 0.654 2.754 0.735 ;
      RECT 2.638 0.312 2.715 0.593 ;
      RECT 2.624 0.312 2.638 0.988 ;
      RECT 2.604 0.538 2.624 0.988 ;
      RECT 2.576 0.538 2.604 1.014 ;
      RECT 2.513 0.933 2.576 1.014 ;
      RECT 2.484 0.189 2.513 0.776 ;
      RECT 2.452 0.189 2.484 0.861 ;
      RECT 2.160 0.414 2.452 0.469 ;
      RECT 2.423 0.695 2.452 0.861 ;
      RECT 2.379 0.806 2.423 0.861 ;
      RECT 2.300 0.524 2.391 0.605 ;
      RECT 2.317 0.806 2.379 1.008 ;
      RECT 1.688 0.954 2.317 1.008 ;
      RECT 2.253 0.550 2.300 0.605 ;
      RECT 2.192 0.550 2.253 0.899 ;
      RECT 1.949 0.844 2.192 0.899 ;
      RECT 2.102 0.279 2.160 0.469 ;
      RECT 2.069 0.279 2.102 0.743 ;
      RECT 2.068 0.292 2.069 0.743 ;
      RECT 2.041 0.414 2.068 0.743 ;
      RECT 2.012 0.662 2.041 0.743 ;
      RECT 1.949 0.193 1.973 0.274 ;
      RECT 1.887 0.193 1.949 0.899 ;
      RECT 1.882 0.193 1.887 0.274 ;
      RECT 1.805 0.542 1.887 0.596 ;
      RECT 1.735 0.369 1.826 0.450 ;
      RECT 1.714 0.529 1.805 0.610 ;
      RECT 1.606 0.382 1.735 0.437 ;
      RECT 1.674 0.900 1.688 1.008 ;
      RECT 1.612 0.885 1.674 1.008 ;
      RECT 1.598 0.885 1.612 0.981 ;
      RECT 1.572 0.189 1.606 0.437 ;
      RECT 1.450 0.885 1.598 0.939 ;
      RECT 1.511 0.189 1.572 0.829 ;
      RECT 1.305 0.189 1.511 0.244 ;
      RECT 1.308 0.995 1.458 1.050 ;
      RECT 1.388 0.419 1.450 0.939 ;
      RECT 1.323 0.419 1.388 0.474 ;
      RECT 1.236 0.790 1.327 0.871 ;
      RECT 1.261 0.331 1.323 0.474 ;
      RECT 1.247 0.933 1.308 1.050 ;
      RECT 0.917 0.933 1.247 0.988 ;
      RECT 0.794 0.817 1.236 0.871 ;
      RECT 1.092 0.179 1.183 0.260 ;
      RECT 0.663 0.193 1.092 0.248 ;
      RECT 0.853 0.320 0.924 0.375 ;
      RECT 0.856 0.933 0.917 1.050 ;
      RECT 0.506 0.995 0.856 1.050 ;
      RECT 0.792 0.302 0.853 0.375 ;
      RECT 0.733 0.817 0.794 0.936 ;
      RECT 0.551 0.302 0.792 0.357 ;
      RECT 0.574 0.881 0.733 0.936 ;
      RECT 0.602 0.154 0.663 0.248 ;
      RECT 0.573 0.724 0.663 0.805 ;
      RECT 0.366 0.154 0.602 0.208 ;
      RECT 0.497 0.724 0.573 0.779 ;
      RECT 0.490 0.302 0.551 0.512 ;
      RECT 0.444 0.858 0.506 1.050 ;
      RECT 0.467 0.692 0.497 0.779 ;
      RECT 0.467 0.457 0.490 0.512 ;
      RECT 0.406 0.457 0.467 0.779 ;
      RECT 0.144 0.858 0.444 0.913 ;
      RECT 0.101 0.713 0.144 0.913 ;
      RECT 0.101 0.340 0.139 0.421 ;
      RECT 0.083 0.340 0.101 0.913 ;
      RECT 0.053 0.340 0.083 0.794 ;
      RECT 0.048 0.340 0.053 0.768 ;
      RECT 0.040 0.354 0.048 0.768 ;
  END
END SDFFNXL

MACRO SDFFNX1
  CLASS CORE ;
  FOREIGN SDFFNX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.762 0.439 0.878 0.567 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.054 0.662 1.069 0.743 ;
      RECT 0.978 0.626 1.054 0.743 ;
      RECT 0.667 0.626 0.978 0.681 ;
      RECT 0.590 0.567 0.667 0.681 ;
      RECT 0.566 0.567 0.590 0.633 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.561 0.283 3.652 0.924 ;
      RECT 3.534 0.843 3.561 0.924 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.405 0.206 3.466 0.814 ;
      RECT 3.385 0.206 3.405 0.306 ;
      RECT 3.169 0.760 3.405 0.814 ;
      RECT 3.278 0.206 3.385 0.261 ;
      RECT 3.187 0.173 3.278 0.261 ;
      RECT 3.078 0.760 3.169 0.840 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.140 0.439 1.176 0.494 ;
      RECT 1.072 0.335 1.140 0.494 ;
      RECT 1.049 0.335 1.072 0.415 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.234 0.525 0.315 0.633 ;
      RECT 0.172 0.512 0.234 0.633 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.497 -0.080 3.700 0.080 ;
      RECT 3.406 -0.080 3.497 0.122 ;
      RECT 3.075 -0.080 3.406 0.080 ;
      RECT 2.985 -0.080 3.075 0.122 ;
      RECT 2.424 -0.080 2.985 0.080 ;
      RECT 2.333 -0.080 2.424 0.359 ;
      RECT 1.791 -0.080 2.333 0.080 ;
      RECT 1.701 -0.080 1.791 0.259 ;
      RECT 0.852 -0.080 1.701 0.080 ;
      RECT 0.761 -0.080 0.852 0.122 ;
      RECT 0.336 -0.080 0.761 0.080 ;
      RECT 0.336 0.335 0.408 0.386 ;
      RECT 0.275 -0.080 0.336 0.386 ;
      RECT 0.000 -0.080 0.275 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.422 1.120 3.700 1.280 ;
      RECT 3.332 1.065 3.422 1.280 ;
      RECT 2.966 1.120 3.332 1.280 ;
      RECT 2.875 1.078 2.966 1.280 ;
      RECT 2.252 1.120 2.875 1.280 ;
      RECT 2.161 1.078 2.252 1.280 ;
      RECT 1.077 1.120 2.161 1.280 ;
      RECT 0.986 1.065 1.077 1.280 ;
      RECT 0.196 1.120 0.986 1.280 ;
      RECT 0.105 1.065 0.196 1.280 ;
      RECT 0.000 1.120 0.105 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.301 0.477 3.340 0.579 ;
      RECT 3.240 0.350 3.301 0.704 ;
      RECT 3.198 0.350 3.240 0.431 ;
      RECT 2.934 0.649 3.240 0.704 ;
      RECT 3.085 0.486 3.175 0.567 ;
      RECT 3.139 0.960 3.169 1.040 ;
      RECT 3.078 0.945 3.139 1.040 ;
      RECT 3.075 0.486 3.085 0.540 ;
      RECT 2.934 0.945 3.078 1.000 ;
      RECT 3.014 0.343 3.075 0.540 ;
      RECT 2.720 0.343 3.014 0.437 ;
      RECT 2.872 0.519 2.934 1.000 ;
      RECT 2.843 0.519 2.872 0.600 ;
      RECT 2.557 0.160 2.867 0.214 ;
      RECT 2.659 0.343 2.720 1.007 ;
      RECT 2.630 0.952 2.659 1.007 ;
      RECT 2.539 0.952 2.630 1.033 ;
      RECT 2.537 0.671 2.597 0.752 ;
      RECT 2.537 0.160 2.557 0.493 ;
      RECT 2.496 0.160 2.537 0.861 ;
      RECT 2.476 0.438 2.496 0.861 ;
      RECT 2.202 0.438 2.476 0.493 ;
      RECT 2.379 0.806 2.476 0.861 ;
      RECT 2.343 0.567 2.404 0.746 ;
      RECT 2.317 0.806 2.379 1.008 ;
      RECT 2.253 0.692 2.343 0.746 ;
      RECT 1.663 0.954 2.317 1.008 ;
      RECT 2.192 0.692 2.253 0.899 ;
      RECT 2.128 0.267 2.202 0.493 ;
      RECT 1.975 0.844 2.192 0.899 ;
      RECT 2.112 0.267 2.128 0.745 ;
      RECT 2.066 0.438 2.112 0.745 ;
      RECT 2.037 0.664 2.066 0.745 ;
      RECT 1.990 0.193 2.005 0.274 ;
      RECT 1.975 0.193 1.990 0.571 ;
      RECT 1.929 0.193 1.975 0.899 ;
      RECT 1.914 0.193 1.929 0.274 ;
      RECT 1.903 0.490 1.929 0.899 ;
      RECT 1.660 0.490 1.903 0.571 ;
      RECT 1.777 0.330 1.867 0.411 ;
      RECT 1.584 0.343 1.777 0.398 ;
      RECT 1.634 0.940 1.663 1.021 ;
      RECT 1.572 0.886 1.634 1.021 ;
      RECT 1.523 0.192 1.584 0.831 ;
      RECT 1.462 0.886 1.572 0.940 ;
      RECT 1.337 0.192 1.523 0.246 ;
      RECT 1.339 0.995 1.478 1.050 ;
      RECT 1.400 0.671 1.462 0.940 ;
      RECT 1.339 0.671 1.400 0.726 ;
      RECT 1.339 0.331 1.353 0.412 ;
      RECT 1.277 0.331 1.339 0.726 ;
      RECT 1.248 0.790 1.339 0.871 ;
      RECT 1.277 0.933 1.339 1.050 ;
      RECT 1.263 0.331 1.277 0.412 ;
      RECT 0.922 0.933 1.277 0.988 ;
      RECT 0.798 0.804 1.248 0.858 ;
      RECT 1.124 0.179 1.215 0.260 ;
      RECT 0.695 0.193 1.124 0.248 ;
      RECT 0.635 0.320 0.960 0.375 ;
      RECT 0.861 0.933 0.922 1.050 ;
      RECT 0.506 0.995 0.861 1.050 ;
      RECT 0.737 0.804 0.798 0.936 ;
      RECT 0.573 0.881 0.737 0.936 ;
      RECT 0.634 0.154 0.695 0.248 ;
      RECT 0.505 0.737 0.675 0.792 ;
      RECT 0.606 0.320 0.635 0.421 ;
      RECT 0.398 0.154 0.634 0.208 ;
      RECT 0.559 0.320 0.606 0.512 ;
      RECT 0.545 0.340 0.559 0.512 ;
      RECT 0.505 0.457 0.545 0.512 ;
      RECT 0.444 0.858 0.506 1.050 ;
      RECT 0.443 0.457 0.505 0.792 ;
      RECT 0.152 0.858 0.444 0.913 ;
      RECT 0.406 0.687 0.443 0.792 ;
      RECT 0.109 0.340 0.200 0.421 ;
      RECT 0.101 0.719 0.152 0.913 ;
      RECT 0.101 0.367 0.109 0.421 ;
      RECT 0.040 0.367 0.101 0.913 ;
  END
END SDFFNX1

MACRO SDFFHQXL
  CLASS CORE ;
  FOREIGN SDFFHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.757 0.439 0.872 0.569 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.960 0.626 1.050 0.717 ;
      RECT 0.663 0.626 0.960 0.681 ;
      RECT 0.586 0.567 0.663 0.681 ;
      RECT 0.562 0.567 0.586 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.443 0.189 3.467 0.839 ;
      RECT 3.406 0.189 3.443 0.894 ;
      RECT 3.382 0.189 3.406 0.244 ;
      RECT 3.382 0.760 3.406 0.894 ;
      RECT 3.333 0.167 3.382 0.244 ;
      RECT 3.110 0.760 3.382 0.840 ;
      RECT 3.243 0.163 3.333 0.244 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.132 0.439 1.168 0.494 ;
      RECT 1.065 0.335 1.132 0.494 ;
      RECT 1.042 0.335 1.065 0.415 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.525 0.313 0.633 ;
      RECT 0.171 0.512 0.232 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.131 -0.080 3.500 0.080 ;
      RECT 3.041 -0.080 3.131 0.122 ;
      RECT 2.374 -0.080 3.041 0.080 ;
      RECT 2.313 -0.080 2.374 0.333 ;
      RECT 1.765 -0.080 2.313 0.080 ;
      RECT 1.704 -0.080 1.765 0.259 ;
      RECT 0.846 -0.080 1.704 0.080 ;
      RECT 0.756 -0.080 0.846 0.122 ;
      RECT 0.334 -0.080 0.756 0.080 ;
      RECT 0.334 0.322 0.419 0.373 ;
      RECT 0.273 -0.080 0.334 0.373 ;
      RECT 0.000 -0.080 0.273 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.988 1.120 3.500 1.280 ;
      RECT 2.898 1.078 2.988 1.280 ;
      RECT 2.237 1.120 2.898 1.280 ;
      RECT 2.146 1.078 2.237 1.280 ;
      RECT 1.151 1.120 2.146 1.280 ;
      RECT 1.061 1.065 1.151 1.280 ;
      RECT 0.292 1.120 1.061 1.280 ;
      RECT 0.202 1.078 0.292 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.332 0.348 3.344 0.429 ;
      RECT 3.271 0.348 3.332 0.705 ;
      RECT 3.253 0.348 3.271 0.429 ;
      RECT 2.991 0.650 3.271 0.705 ;
      RECT 3.131 0.486 3.210 0.567 ;
      RECT 3.100 0.954 3.190 1.048 ;
      RECT 3.070 0.382 3.131 0.567 ;
      RECT 2.991 0.954 3.100 1.008 ;
      RECT 2.809 0.382 3.070 0.437 ;
      RECT 2.930 0.519 2.991 1.008 ;
      RECT 2.901 0.519 2.930 0.600 ;
      RECT 2.496 0.208 2.925 0.263 ;
      RECT 2.748 0.326 2.809 1.010 ;
      RECT 2.665 0.955 2.748 1.010 ;
      RECT 2.626 0.318 2.687 0.874 ;
      RECT 2.575 0.955 2.665 1.036 ;
      RECT 2.557 0.318 2.626 0.399 ;
      RECT 2.459 0.819 2.626 0.874 ;
      RECT 2.504 0.454 2.565 0.760 ;
      RECT 2.496 0.454 2.504 0.508 ;
      RECT 2.327 0.705 2.504 0.760 ;
      RECT 2.435 0.208 2.496 0.508 ;
      RECT 2.398 0.819 2.459 0.996 ;
      RECT 2.266 0.454 2.435 0.508 ;
      RECT 2.312 0.567 2.402 0.648 ;
      RECT 2.266 0.705 2.327 1.008 ;
      RECT 2.205 0.593 2.312 0.648 ;
      RECT 2.205 0.420 2.266 0.508 ;
      RECT 1.655 0.954 2.266 1.008 ;
      RECT 2.174 0.420 2.205 0.475 ;
      RECT 2.144 0.593 2.205 0.899 ;
      RECT 2.123 0.279 2.177 0.360 ;
      RECT 1.926 0.844 2.144 0.899 ;
      RECT 2.099 0.150 2.123 0.360 ;
      RECT 2.083 0.150 2.099 0.385 ;
      RECT 2.062 0.150 2.083 0.745 ;
      RECT 2.038 0.292 2.062 0.745 ;
      RECT 2.022 0.330 2.038 0.745 ;
      RECT 1.926 0.193 1.977 0.275 ;
      RECT 1.916 0.193 1.926 0.899 ;
      RECT 1.865 0.220 1.916 0.899 ;
      RECT 1.739 0.533 1.865 0.588 ;
      RECT 1.743 0.346 1.804 0.429 ;
      RECT 1.574 0.346 1.743 0.401 ;
      RECT 1.649 0.507 1.739 0.588 ;
      RECT 1.652 0.933 1.655 1.008 ;
      RECT 1.562 0.933 1.652 1.021 ;
      RECT 1.513 0.192 1.574 0.876 ;
      RECT 1.452 0.933 1.562 0.988 ;
      RECT 1.328 0.192 1.513 0.246 ;
      RECT 1.391 0.671 1.452 0.988 ;
      RECT 1.344 0.671 1.391 0.726 ;
      RECT 1.000 0.933 1.391 0.988 ;
      RECT 1.283 0.331 1.344 0.726 ;
      RECT 1.240 0.790 1.330 0.871 ;
      RECT 1.254 0.331 1.283 0.412 ;
      RECT 0.878 0.817 1.240 0.871 ;
      RECT 1.116 0.179 1.206 0.260 ;
      RECT 0.691 0.193 1.116 0.248 ;
      RECT 0.939 0.933 1.000 1.050 ;
      RECT 0.631 0.323 0.953 0.377 ;
      RECT 0.502 0.995 0.939 1.050 ;
      RECT 0.817 0.817 0.878 0.936 ;
      RECT 0.569 0.881 0.817 0.936 ;
      RECT 0.501 0.737 0.756 0.792 ;
      RECT 0.630 0.154 0.691 0.248 ;
      RECT 0.602 0.323 0.631 0.417 ;
      RECT 0.395 0.154 0.630 0.208 ;
      RECT 0.541 0.323 0.602 0.511 ;
      RECT 0.501 0.456 0.541 0.511 ;
      RECT 0.441 0.858 0.502 1.050 ;
      RECT 0.440 0.456 0.501 0.792 ;
      RECT 0.151 0.858 0.441 0.913 ;
      RECT 0.403 0.687 0.440 0.768 ;
      RECT 0.109 0.336 0.199 0.417 ;
      RECT 0.101 0.719 0.151 0.913 ;
      RECT 0.101 0.362 0.109 0.417 ;
      RECT 0.040 0.362 0.101 0.913 ;
  END
END SDFFHQXL

MACRO SDFFHQX4
  CLASS CORE ;
  FOREIGN SDFFHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.839 0.433 0.871 0.533 ;
      RECT 0.750 0.433 0.839 0.546 ;
      RECT 0.729 0.433 0.750 0.500 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.926 0.593 1.015 0.674 ;
      RECT 0.690 0.601 0.926 0.656 ;
      RECT 0.629 0.567 0.690 0.656 ;
      RECT 0.527 0.567 0.629 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.282 0.433 4.290 0.767 ;
      RECT 4.193 0.325 4.282 0.767 ;
      RECT 4.191 0.433 4.193 0.767 ;
      RECT 4.130 0.671 4.191 0.752 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.150 0.356 1.156 0.439 ;
      RECT 1.150 0.573 1.155 0.627 ;
      RECT 1.088 0.356 1.150 0.627 ;
      RECT 1.067 0.356 1.088 0.437 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.152 0.524 0.290 0.627 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.450 -0.080 4.500 0.080 ;
      RECT 4.361 -0.080 4.450 0.215 ;
      RECT 4.115 -0.080 4.361 0.080 ;
      RECT 4.025 -0.080 4.115 0.212 ;
      RECT 3.721 -0.080 4.025 0.080 ;
      RECT 3.632 -0.080 3.721 0.122 ;
      RECT 3.245 -0.080 3.632 0.080 ;
      RECT 3.185 -0.080 3.245 0.287 ;
      RECT 2.422 -0.080 3.185 0.080 ;
      RECT 2.361 -0.080 2.422 0.311 ;
      RECT 1.767 -0.080 2.361 0.080 ;
      RECT 1.678 -0.080 1.767 0.287 ;
      RECT 0.844 -0.080 1.678 0.080 ;
      RECT 0.755 -0.080 0.844 0.122 ;
      RECT 0.338 -0.080 0.755 0.080 ;
      RECT 0.338 0.359 0.346 0.410 ;
      RECT 0.249 -0.080 0.338 0.410 ;
      RECT 0.000 -0.080 0.249 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.389 1.120 4.500 1.280 ;
      RECT 4.299 0.989 4.389 1.280 ;
      RECT 4.040 1.120 4.299 1.280 ;
      RECT 3.951 1.078 4.040 1.280 ;
      RECT 3.687 1.120 3.951 1.280 ;
      RECT 3.060 1.078 3.687 1.280 ;
      RECT 2.373 1.120 3.060 1.280 ;
      RECT 2.284 1.078 2.373 1.280 ;
      RECT 1.479 1.120 2.284 1.280 ;
      RECT 1.390 1.078 1.479 1.280 ;
      RECT 0.337 1.120 1.390 1.280 ;
      RECT 0.248 1.078 0.337 1.280 ;
      RECT 0.000 1.120 0.248 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.923 0.264 3.931 0.345 ;
      RECT 3.863 0.264 3.923 0.907 ;
      RECT 3.842 0.264 3.863 0.571 ;
      RECT 3.799 0.826 3.863 0.907 ;
      RECT 3.699 0.490 3.842 0.571 ;
      RECT 3.636 0.650 3.802 0.731 ;
      RECT 3.576 0.357 3.636 0.886 ;
      RECT 3.469 0.357 3.576 0.412 ;
      RECT 3.363 0.831 3.576 0.886 ;
      RECT 3.414 0.467 3.475 0.768 ;
      RECT 3.380 0.150 3.469 0.412 ;
      RECT 3.003 0.467 3.414 0.521 ;
      RECT 3.241 0.713 3.414 0.768 ;
      RECT 3.125 0.357 3.380 0.412 ;
      RECT 3.303 0.831 3.363 1.008 ;
      RECT 3.265 0.577 3.354 0.658 ;
      RECT 2.761 0.954 3.303 1.008 ;
      RECT 3.121 0.604 3.265 0.658 ;
      RECT 3.181 0.713 3.241 0.898 ;
      RECT 2.573 0.843 3.181 0.898 ;
      RECT 3.064 0.223 3.125 0.412 ;
      RECT 3.060 0.604 3.121 0.787 ;
      RECT 2.814 0.223 3.064 0.277 ;
      RECT 2.685 0.732 3.060 0.787 ;
      RECT 2.942 0.348 3.003 0.521 ;
      RECT 2.911 0.596 3.000 0.677 ;
      RECT 2.913 0.348 2.942 0.429 ;
      RECT 2.628 0.374 2.913 0.429 ;
      RECT 2.807 0.598 2.911 0.652 ;
      RECT 2.725 0.223 2.814 0.304 ;
      RECT 2.747 0.490 2.807 0.652 ;
      RECT 2.672 0.954 2.761 1.035 ;
      RECT 2.510 0.490 2.747 0.545 ;
      RECT 2.596 0.605 2.685 0.787 ;
      RECT 2.567 0.245 2.628 0.429 ;
      RECT 2.347 0.732 2.596 0.787 ;
      RECT 2.483 0.843 2.573 0.924 ;
      RECT 2.536 0.245 2.567 0.326 ;
      RECT 2.481 0.490 2.510 0.571 ;
      RECT 2.420 0.381 2.481 0.571 ;
      RECT 2.301 0.381 2.420 0.436 ;
      RECT 2.310 0.530 2.347 0.993 ;
      RECT 2.287 0.504 2.310 0.993 ;
      RECT 2.241 0.158 2.301 0.436 ;
      RECT 2.221 0.504 2.287 0.585 ;
      RECT 1.634 0.938 2.287 0.993 ;
      RECT 1.956 0.158 2.241 0.213 ;
      RECT 2.198 0.789 2.226 0.870 ;
      RECT 2.161 0.679 2.198 0.870 ;
      RECT 2.161 0.269 2.181 0.402 ;
      RECT 2.137 0.269 2.161 0.870 ;
      RECT 2.120 0.269 2.137 0.733 ;
      RECT 2.101 0.348 2.120 0.733 ;
      RECT 2.010 0.454 2.101 0.535 ;
      RECT 1.952 0.790 2.042 0.871 ;
      RECT 1.950 0.158 1.956 0.354 ;
      RECT 1.950 0.790 1.952 0.858 ;
      RECT 1.896 0.158 1.950 0.858 ;
      RECT 1.889 0.273 1.896 0.858 ;
      RECT 1.867 0.273 1.889 0.354 ;
      RECT 1.689 0.612 1.889 0.693 ;
      RECT 1.740 0.450 1.829 0.531 ;
      RECT 1.524 0.450 1.740 0.505 ;
      RECT 1.545 0.938 1.634 1.019 ;
      RECT 1.403 0.939 1.545 0.994 ;
      RECT 1.463 0.163 1.524 0.855 ;
      RECT 1.322 0.163 1.463 0.218 ;
      RECT 1.343 0.357 1.403 0.994 ;
      RECT 1.337 0.357 1.343 0.412 ;
      RECT 1.145 0.939 1.343 0.994 ;
      RECT 1.248 0.331 1.337 0.412 ;
      RECT 1.193 0.776 1.282 0.857 ;
      RECT 1.112 0.160 1.201 0.246 ;
      RECT 1.012 0.802 1.193 0.857 ;
      RECT 1.084 0.939 1.145 1.050 ;
      RECT 0.490 0.192 1.112 0.246 ;
      RECT 0.483 0.995 1.084 1.050 ;
      RECT 0.952 0.802 1.012 0.936 ;
      RECT 0.580 0.318 0.952 0.373 ;
      RECT 0.543 0.881 0.952 0.936 ;
      RECT 0.606 0.724 0.695 0.805 ;
      RECT 0.509 0.724 0.606 0.779 ;
      RECT 0.551 0.318 0.580 0.425 ;
      RECT 0.490 0.318 0.551 0.512 ;
      RECT 0.467 0.692 0.509 0.779 ;
      RECT 0.399 0.154 0.490 0.246 ;
      RECT 0.467 0.457 0.490 0.512 ;
      RECT 0.422 0.877 0.483 1.050 ;
      RECT 0.406 0.457 0.467 0.779 ;
      RECT 0.136 0.877 0.422 0.932 ;
      RECT 0.092 0.344 0.157 0.425 ;
      RECT 0.122 0.739 0.136 0.932 ;
      RECT 0.092 0.688 0.122 0.932 ;
      RECT 0.068 0.344 0.092 0.932 ;
      RECT 0.047 0.369 0.068 0.932 ;
      RECT 0.031 0.369 0.047 0.743 ;
  END
END SDFFHQX4

MACRO SDFFHQX1
  CLASS CORE ;
  FOREIGN SDFFHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.737 0.433 0.924 0.548 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.960 0.614 1.050 0.743 ;
      RECT 0.663 0.614 0.960 0.669 ;
      RECT 0.563 0.567 0.663 0.669 ;
      RECT 0.562 0.567 0.563 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.443 0.188 3.467 0.839 ;
      RECT 3.406 0.188 3.443 0.894 ;
      RECT 3.382 0.188 3.406 0.243 ;
      RECT 3.382 0.760 3.406 0.894 ;
      RECT 3.333 0.167 3.382 0.243 ;
      RECT 3.100 0.760 3.382 0.840 ;
      RECT 3.243 0.162 3.333 0.243 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.132 0.439 1.168 0.494 ;
      RECT 1.065 0.335 1.132 0.494 ;
      RECT 1.042 0.335 1.065 0.415 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.525 0.313 0.633 ;
      RECT 0.171 0.512 0.232 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.131 -0.080 3.500 0.080 ;
      RECT 3.041 -0.080 3.131 0.122 ;
      RECT 2.374 -0.080 3.041 0.080 ;
      RECT 2.313 -0.080 2.374 0.333 ;
      RECT 1.779 -0.080 2.313 0.080 ;
      RECT 1.689 -0.080 1.779 0.259 ;
      RECT 0.846 -0.080 1.689 0.080 ;
      RECT 0.756 -0.080 0.846 0.122 ;
      RECT 0.334 -0.080 0.756 0.080 ;
      RECT 0.334 0.322 0.406 0.373 ;
      RECT 0.273 -0.080 0.334 0.373 ;
      RECT 0.000 -0.080 0.273 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.391 1.120 3.500 1.280 ;
      RECT 3.301 1.065 3.391 1.280 ;
      RECT 2.988 1.120 3.301 1.280 ;
      RECT 2.898 1.078 2.988 1.280 ;
      RECT 2.211 1.120 2.898 1.280 ;
      RECT 1.872 1.078 2.211 1.280 ;
      RECT 1.151 1.120 1.872 1.280 ;
      RECT 1.061 1.065 1.151 1.280 ;
      RECT 0.292 1.120 1.061 1.280 ;
      RECT 0.202 1.078 0.292 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.283 0.348 3.344 0.705 ;
      RECT 3.253 0.348 3.283 0.429 ;
      RECT 2.991 0.650 3.283 0.705 ;
      RECT 3.149 0.486 3.210 0.567 ;
      RECT 3.110 0.980 3.190 1.035 ;
      RECT 3.131 0.486 3.149 0.540 ;
      RECT 3.070 0.382 3.131 0.540 ;
      RECT 3.049 0.954 3.110 1.035 ;
      RECT 2.809 0.382 3.070 0.437 ;
      RECT 2.991 0.954 3.049 1.008 ;
      RECT 2.930 0.519 2.991 1.008 ;
      RECT 2.901 0.519 2.930 0.600 ;
      RECT 2.834 0.195 2.925 0.276 ;
      RECT 2.496 0.208 2.834 0.263 ;
      RECT 2.748 0.343 2.809 1.008 ;
      RECT 2.654 0.954 2.748 1.008 ;
      RECT 2.626 0.344 2.687 0.883 ;
      RECT 2.564 0.954 2.654 1.035 ;
      RECT 2.618 0.344 2.626 0.399 ;
      RECT 2.449 0.829 2.626 0.883 ;
      RECT 2.557 0.318 2.618 0.399 ;
      RECT 2.520 0.671 2.565 0.770 ;
      RECT 2.496 0.455 2.520 0.770 ;
      RECT 2.459 0.208 2.496 0.770 ;
      RECT 2.435 0.208 2.459 0.510 ;
      RECT 2.327 0.715 2.459 0.770 ;
      RECT 2.388 0.829 2.449 0.996 ;
      RECT 2.174 0.420 2.435 0.475 ;
      RECT 2.205 0.567 2.388 0.651 ;
      RECT 2.266 0.715 2.327 1.008 ;
      RECT 1.652 0.954 2.266 1.008 ;
      RECT 2.144 0.567 2.205 0.899 ;
      RECT 2.137 0.279 2.177 0.360 ;
      RECT 1.941 0.844 2.144 0.899 ;
      RECT 2.108 0.150 2.137 0.360 ;
      RECT 2.083 0.150 2.108 0.385 ;
      RECT 2.047 0.150 2.083 0.745 ;
      RECT 2.022 0.330 2.047 0.745 ;
      RECT 1.941 0.193 1.977 0.275 ;
      RECT 1.916 0.193 1.941 0.899 ;
      RECT 1.880 0.220 1.916 0.899 ;
      RECT 1.710 0.507 1.880 0.588 ;
      RECT 1.729 0.348 1.819 0.429 ;
      RECT 1.574 0.374 1.729 0.429 ;
      RECT 1.562 0.940 1.652 1.021 ;
      RECT 1.513 0.192 1.574 0.876 ;
      RECT 1.452 0.940 1.562 0.995 ;
      RECT 1.419 0.192 1.513 0.260 ;
      RECT 1.391 0.357 1.452 0.995 ;
      RECT 1.328 0.179 1.419 0.260 ;
      RECT 1.344 0.357 1.391 0.412 ;
      RECT 1.000 0.940 1.391 0.995 ;
      RECT 1.254 0.331 1.344 0.412 ;
      RECT 1.240 0.790 1.330 0.871 ;
      RECT 0.878 0.817 1.240 0.871 ;
      RECT 1.116 0.179 1.206 0.260 ;
      RECT 0.691 0.205 1.116 0.260 ;
      RECT 0.939 0.940 1.000 1.050 ;
      RECT 0.631 0.320 0.953 0.375 ;
      RECT 0.502 0.995 0.939 1.050 ;
      RECT 0.817 0.817 0.878 0.936 ;
      RECT 0.569 0.881 0.817 0.936 ;
      RECT 0.634 0.724 0.724 0.805 ;
      RECT 0.630 0.154 0.691 0.260 ;
      RECT 0.501 0.724 0.634 0.779 ;
      RECT 0.541 0.320 0.631 0.421 ;
      RECT 0.395 0.154 0.630 0.208 ;
      RECT 0.528 0.367 0.541 0.421 ;
      RECT 0.501 0.367 0.528 0.511 ;
      RECT 0.441 0.858 0.502 1.050 ;
      RECT 0.467 0.367 0.501 0.779 ;
      RECT 0.440 0.456 0.467 0.779 ;
      RECT 0.151 0.858 0.441 0.913 ;
      RECT 0.403 0.687 0.440 0.779 ;
      RECT 0.109 0.340 0.199 0.421 ;
      RECT 0.101 0.719 0.151 0.913 ;
      RECT 0.101 0.367 0.109 0.421 ;
      RECT 0.040 0.367 0.101 0.913 ;
  END
END SDFFHQX1

MACRO SDFFXL
  CLASS CORE ;
  FOREIGN SDFFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.715 0.433 0.838 0.500 ;
      RECT 0.627 0.412 0.715 0.500 ;
      RECT 0.613 0.412 0.627 0.467 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.947 0.619 1.037 0.700 ;
      RECT 0.843 0.619 0.947 0.674 ;
      RECT 0.782 0.567 0.843 0.674 ;
      RECT 0.587 0.567 0.782 0.633 ;
      RECT 0.497 0.558 0.587 0.639 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.443 0.837 3.452 0.918 ;
      RECT 3.399 0.282 3.443 0.918 ;
      RECT 3.382 0.260 3.399 0.918 ;
      RECT 3.309 0.260 3.382 0.340 ;
      RECT 3.362 0.837 3.382 0.918 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.175 0.163 3.177 0.248 ;
      RECT 3.085 0.150 3.175 0.248 ;
      RECT 3.090 0.513 3.139 0.819 ;
      RECT 3.078 0.513 3.090 0.845 ;
      RECT 3.021 0.193 3.085 0.248 ;
      RECT 3.021 0.513 3.078 0.568 ;
      RECT 3.000 0.764 3.078 0.845 ;
      RECT 2.960 0.193 3.021 0.568 ;
      RECT 2.857 0.300 2.960 0.367 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.010 0.314 1.100 0.494 ;
      RECT 0.932 0.439 1.010 0.494 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.537 0.313 0.633 ;
      RECT 0.212 0.524 0.232 0.633 ;
      RECT 0.171 0.524 0.212 0.632 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.389 -0.080 3.500 0.080 ;
      RECT 3.298 -0.080 3.389 0.122 ;
      RECT 2.974 -0.080 3.298 0.080 ;
      RECT 2.884 -0.080 2.974 0.122 ;
      RECT 2.327 -0.080 2.884 0.080 ;
      RECT 2.237 -0.080 2.327 0.345 ;
      RECT 1.716 -0.080 2.237 0.080 ;
      RECT 1.625 -0.080 1.716 0.259 ;
      RECT 0.814 -0.080 1.625 0.080 ;
      RECT 0.724 -0.080 0.814 0.122 ;
      RECT 0.302 -0.080 0.724 0.080 ;
      RECT 0.302 0.322 0.350 0.373 ;
      RECT 0.260 -0.080 0.302 0.373 ;
      RECT 0.241 -0.080 0.260 0.360 ;
      RECT 0.000 -0.080 0.241 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.265 1.120 3.500 1.280 ;
      RECT 3.175 1.065 3.265 1.280 ;
      RECT 2.877 1.120 3.175 1.280 ;
      RECT 2.787 1.078 2.877 1.280 ;
      RECT 2.218 1.120 2.787 1.280 ;
      RECT 1.879 1.078 2.218 1.280 ;
      RECT 1.066 1.120 1.879 1.280 ;
      RECT 0.976 1.065 1.066 1.280 ;
      RECT 0.292 1.120 0.976 1.280 ;
      RECT 0.202 1.078 0.292 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.240 0.401 3.301 0.995 ;
      RECT 3.171 0.401 3.240 0.456 ;
      RECT 3.112 0.940 3.240 0.995 ;
      RECT 3.110 0.324 3.171 0.456 ;
      RECT 3.051 0.940 3.112 1.036 ;
      RECT 2.980 0.954 3.051 1.036 ;
      RECT 2.926 0.623 3.016 0.704 ;
      RECT 2.763 0.954 2.980 1.008 ;
      RECT 2.885 0.623 2.926 0.677 ;
      RECT 2.824 0.438 2.885 0.677 ;
      RECT 2.666 0.438 2.824 0.493 ;
      RECT 2.702 0.596 2.763 1.008 ;
      RECT 2.465 0.160 2.740 0.214 ;
      RECT 2.637 0.302 2.666 0.493 ;
      RECT 2.576 0.302 2.637 0.988 ;
      RECT 2.568 0.933 2.576 0.988 ;
      RECT 2.478 0.933 2.568 1.014 ;
      RECT 2.465 0.695 2.470 0.776 ;
      RECT 2.441 0.160 2.465 0.776 ;
      RECT 2.417 0.160 2.441 0.856 ;
      RECT 2.404 0.160 2.417 1.008 ;
      RECT 2.157 0.414 2.404 0.469 ;
      RECT 2.380 0.695 2.404 1.008 ;
      RECT 2.356 0.801 2.380 1.008 ;
      RECT 1.643 0.954 2.356 1.008 ;
      RECT 2.282 0.524 2.341 0.606 ;
      RECT 2.238 0.524 2.282 0.746 ;
      RECT 2.221 0.524 2.238 0.899 ;
      RECT 2.177 0.692 2.221 0.899 ;
      RECT 1.835 0.844 2.177 0.899 ;
      RECT 2.096 0.414 2.157 0.598 ;
      RECT 2.088 0.279 2.115 0.360 ;
      RECT 2.035 0.150 2.088 0.360 ;
      RECT 2.035 0.662 2.060 0.743 ;
      RECT 1.974 0.150 2.035 0.743 ;
      RECT 1.970 0.662 1.974 0.743 ;
      RECT 1.852 0.193 1.913 0.577 ;
      RECT 1.835 0.523 1.852 0.577 ;
      RECT 1.774 0.523 1.835 0.899 ;
      RECT 1.700 0.379 1.790 0.460 ;
      RECT 1.673 0.571 1.774 0.652 ;
      RECT 1.562 0.379 1.700 0.433 ;
      RECT 1.552 0.940 1.643 1.021 ;
      RECT 1.537 0.202 1.562 0.433 ;
      RECT 1.415 0.940 1.552 0.995 ;
      RECT 1.476 0.202 1.537 0.876 ;
      RECT 1.355 0.202 1.476 0.257 ;
      RECT 1.354 0.671 1.415 0.995 ;
      RECT 1.265 0.176 1.355 0.257 ;
      RECT 1.263 0.671 1.354 0.726 ;
      RECT 0.915 0.940 1.354 0.995 ;
      RECT 1.202 0.790 1.293 0.871 ;
      RECT 1.202 0.331 1.263 0.726 ;
      RECT 0.793 0.804 1.202 0.858 ;
      RECT 1.074 0.179 1.164 0.260 ;
      RECT 0.659 0.193 1.074 0.248 ;
      RECT 0.854 0.940 0.915 1.050 ;
      RECT 0.785 0.302 0.888 0.375 ;
      RECT 0.459 0.995 0.854 1.050 ;
      RECT 0.732 0.804 0.793 0.936 ;
      RECT 0.548 0.302 0.785 0.357 ;
      RECT 0.555 0.881 0.732 0.936 ;
      RECT 0.598 0.154 0.659 0.248 ;
      RECT 0.566 0.726 0.656 0.821 ;
      RECT 0.363 0.154 0.598 0.208 ;
      RECT 0.493 0.726 0.566 0.781 ;
      RECT 0.487 0.302 0.548 0.499 ;
      RECT 0.436 0.700 0.493 0.781 ;
      RECT 0.436 0.444 0.487 0.499 ;
      RECT 0.398 0.937 0.459 1.050 ;
      RECT 0.375 0.444 0.436 0.781 ;
      RECT 0.143 0.937 0.398 0.992 ;
      RECT 0.101 0.718 0.143 0.992 ;
      RECT 0.101 0.340 0.138 0.421 ;
      RECT 0.082 0.340 0.101 0.992 ;
      RECT 0.040 0.340 0.082 0.800 ;
  END
END SDFFXL

MACRO OR4X2
  CLASS CORE ;
  FOREIGN OR4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.997 0.182 1.061 1.010 ;
      RECT 0.942 0.182 0.997 0.375 ;
      RECT 0.953 0.700 0.997 1.010 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.728 0.700 0.878 0.767 ;
      RECT 0.664 0.552 0.728 0.767 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.406 0.527 0.556 0.633 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.167 0.364 0.264 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.433 0.151 0.567 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.646 -0.080 1.100 0.080 ;
      RECT 0.551 -0.080 0.646 0.122 ;
      RECT 0.144 -0.080 0.551 0.080 ;
      RECT 0.050 -0.080 0.144 0.122 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.836 1.120 1.100 1.280 ;
      RECT 0.742 1.078 0.836 1.280 ;
      RECT 0.000 1.120 0.742 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.876 0.462 0.918 0.576 ;
      RECT 0.812 0.333 0.876 0.576 ;
      RECT 0.669 0.333 0.812 0.388 ;
      RECT 0.575 0.320 0.669 0.401 ;
      RECT 0.285 0.333 0.575 0.388 ;
      RECT 0.279 0.320 0.285 0.388 ;
      RECT 0.215 0.320 0.279 0.717 ;
      RECT 0.144 0.662 0.215 0.717 ;
      RECT 0.081 0.662 0.144 0.924 ;
      RECT 0.050 0.731 0.081 0.924 ;
  END
END OR4X2

MACRO OR4X1
  CLASS CORE ;
  FOREIGN OR4X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.056 0.833 1.061 0.921 ;
      RECT 0.992 0.226 1.056 0.921 ;
      RECT 0.950 0.226 0.992 0.307 ;
      RECT 0.900 0.833 0.992 0.921 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.754 0.555 0.886 0.665 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.486 0.555 0.550 0.767 ;
      RECT 0.406 0.693 0.486 0.767 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.517 0.356 0.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.656 0.156 0.773 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.833 -0.080 1.100 0.080 ;
      RECT 0.739 -0.080 0.833 0.122 ;
      RECT 0.311 -0.080 0.739 0.080 ;
      RECT 0.217 -0.080 0.311 0.122 ;
      RECT 0.000 -0.080 0.217 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.783 1.120 1.100 1.280 ;
      RECT 0.689 1.078 0.783 1.280 ;
      RECT 0.000 1.120 0.689 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.689 0.394 0.915 0.477 ;
      RECT 0.625 0.281 0.689 0.932 ;
      RECT 0.572 0.281 0.625 0.362 ;
      RECT 0.150 0.877 0.625 0.932 ;
      RECT 0.222 0.281 0.572 0.336 ;
      RECT 0.158 0.281 0.222 0.424 ;
      RECT 0.128 0.343 0.158 0.424 ;
      RECT 0.056 0.864 0.150 0.945 ;
  END
END OR4X1

MACRO OR3XL
  CLASS CORE ;
  FOREIGN OR3XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.791 0.348 0.854 0.871 ;
      RECT 0.749 0.348 0.791 0.429 ;
      RECT 0.758 0.706 0.791 0.871 ;
      RECT 0.715 0.790 0.758 0.871 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.637 0.545 0.767 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.433 0.402 0.556 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.206 0.636 0.269 1.027 ;
      RECT 0.164 0.636 0.206 0.721 ;
      RECT 0.059 0.973 0.206 1.027 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.687 -0.080 0.900 0.080 ;
      RECT 0.595 -0.080 0.687 0.122 ;
      RECT 0.153 -0.080 0.595 0.080 ;
      RECT 0.060 -0.080 0.153 0.122 ;
      RECT 0.000 -0.080 0.060 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.655 1.120 0.900 1.280 ;
      RECT 0.562 1.078 0.655 1.280 ;
      RECT 0.000 1.120 0.562 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.635 0.498 0.728 0.579 ;
      RECT 0.627 0.498 0.635 0.552 ;
      RECT 0.565 0.294 0.627 0.552 ;
      RECT 0.496 0.294 0.565 0.349 ;
      RECT 0.404 0.192 0.496 0.349 ;
      RECT 0.142 0.294 0.404 0.349 ;
      RECT 0.101 0.294 0.142 0.429 ;
      RECT 0.101 0.777 0.142 0.858 ;
      RECT 0.038 0.294 0.101 0.858 ;
  END
END OR3XL

MACRO OR3X4
  CLASS CORE ;
  FOREIGN OR3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.207 0.679 1.339 0.767 ;
      RECT 1.207 0.331 1.274 0.412 ;
      RECT 1.104 0.331 1.207 0.767 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.917 0.413 0.966 0.468 ;
      RECT 0.855 0.413 0.917 0.758 ;
      RECT 0.831 0.700 0.855 0.758 ;
      RECT 0.769 0.704 0.831 0.758 ;
      RECT 0.696 0.704 0.769 0.767 ;
      RECT 0.634 0.704 0.696 0.804 ;
      RECT 0.236 0.749 0.634 0.804 ;
      RECT 0.215 0.700 0.236 0.804 ;
      RECT 0.154 0.604 0.215 0.804 ;
      RECT 0.124 0.604 0.154 0.775 ;
      RECT 0.038 0.681 0.124 0.775 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.667 0.457 0.758 0.583 ;
      RECT 0.298 0.457 0.667 0.512 ;
      RECT 0.264 0.439 0.298 0.512 ;
      RECT 0.172 0.431 0.264 0.512 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.392 0.567 0.548 0.694 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.495 -0.080 1.600 0.080 ;
      RECT 1.403 -0.080 1.495 0.122 ;
      RECT 1.049 -0.080 1.403 0.080 ;
      RECT 0.958 -0.080 1.049 0.122 ;
      RECT 0.621 -0.080 0.958 0.080 ;
      RECT 0.529 -0.080 0.621 0.222 ;
      RECT 0.000 -0.080 0.529 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.510 1.120 1.600 1.280 ;
      RECT 1.418 0.983 1.510 1.280 ;
      RECT 1.153 1.120 1.418 1.280 ;
      RECT 1.061 0.983 1.153 1.280 ;
      RECT 0.140 1.120 1.061 1.280 ;
      RECT 0.048 1.078 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.401 0.213 1.463 0.898 ;
      RECT 0.835 0.213 1.401 0.268 ;
      RECT 1.332 0.532 1.401 0.613 ;
      RECT 0.853 0.843 1.401 0.898 ;
      RECT 0.791 0.843 0.853 0.951 ;
      RECT 0.831 0.213 0.835 0.358 ;
      RECT 0.739 0.162 0.831 0.358 ;
      RECT 0.646 0.896 0.791 0.951 ;
      RECT 0.413 0.304 0.739 0.358 ;
      RECT 0.555 0.896 0.646 0.977 ;
      RECT 0.322 0.162 0.413 0.358 ;
  END
END OR3X4

MACRO OR2X4
  CLASS CORE ;
  FOREIGN OR2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.694 0.324 0.733 0.405 ;
      RECT 0.696 0.652 0.700 0.733 ;
      RECT 0.694 0.624 0.696 0.733 ;
      RECT 0.606 0.300 0.694 0.733 ;
      RECT 0.589 0.300 0.606 0.633 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.343 0.479 0.511 0.663 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.392 0.144 0.556 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.922 -0.080 1.100 0.080 ;
      RECT 0.828 -0.080 0.922 0.122 ;
      RECT 0.556 -0.080 0.828 0.080 ;
      RECT 0.461 -0.080 0.556 0.214 ;
      RECT 0.144 -0.080 0.461 0.080 ;
      RECT 0.050 -0.080 0.144 0.290 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.889 1.120 1.100 1.280 ;
      RECT 0.794 1.078 0.889 1.280 ;
      RECT 0.511 1.120 0.794 1.280 ;
      RECT 0.417 1.078 0.511 1.280 ;
      RECT 0.000 1.120 0.417 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.836 0.500 0.867 0.581 ;
      RECT 0.772 0.500 0.836 0.843 ;
      RECT 0.278 0.788 0.772 0.843 ;
      RECT 0.278 0.276 0.344 0.357 ;
      RECT 0.214 0.276 0.278 0.843 ;
      RECT 0.050 0.669 0.214 0.750 ;
  END
END OR2X4

MACRO OR2X2
  CLASS CORE ;
  FOREIGN OR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.589 0.196 0.650 0.914 ;
      RECT 0.548 0.196 0.589 0.389 ;
      RECT 0.546 0.721 0.589 0.914 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.414 0.337 0.558 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.393 0.138 0.544 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 -0.080 0.700 0.080 ;
      RECT 0.345 -0.080 0.435 0.122 ;
      RECT 0.138 -0.080 0.345 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 1.120 0.700 1.280 ;
      RECT 0.345 1.078 0.435 1.280 ;
      RECT 0.000 1.120 0.345 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.460 0.502 0.528 0.583 ;
      RECT 0.399 0.279 0.460 0.776 ;
      RECT 0.286 0.279 0.399 0.333 ;
      RECT 0.138 0.721 0.399 0.776 ;
      RECT 0.196 0.252 0.286 0.333 ;
      RECT 0.048 0.721 0.138 0.802 ;
  END
END OR2X2

MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.597 0.314 0.658 0.867 ;
      RECT 0.562 0.314 0.597 0.395 ;
      RECT 0.562 0.695 0.597 0.867 ;
      RECT 0.553 0.786 0.562 0.867 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 0.567 0.323 0.767 ;
      RECT 0.228 0.567 0.313 0.771 ;
      RECT 0.212 0.700 0.228 0.771 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.474 0.154 0.638 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.369 -0.080 0.700 0.080 ;
      RECT 0.119 -0.080 0.369 0.122 ;
      RECT 0.000 -0.080 0.119 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.384 1.120 0.700 1.280 ;
      RECT 0.290 1.059 0.384 1.280 ;
      RECT 0.000 1.120 0.290 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.471 0.512 0.536 0.593 ;
      RECT 0.410 0.313 0.471 0.906 ;
      RECT 0.215 0.313 0.410 0.368 ;
      RECT 0.143 0.851 0.410 0.906 ;
      RECT 0.118 0.313 0.215 0.405 ;
      RECT 0.053 0.838 0.143 0.919 ;
  END
END OR2X1

MACRO OAI33X1
  CLASS CORE ;
  FOREIGN OAI33X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.310 0.573 1.343 0.627 ;
      RECT 1.249 0.268 1.310 0.887 ;
      RECT 1.193 0.268 1.249 0.414 ;
      RECT 0.626 0.832 1.249 0.887 ;
      RECT 0.902 0.360 1.193 0.414 ;
      RECT 0.811 0.313 0.902 0.414 ;
      RECT 0.536 0.819 0.626 0.900 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.464 0.141 0.633 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.469 0.379 0.633 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.541 0.537 0.570 0.618 ;
      RECT 0.480 0.537 0.541 0.761 ;
      RECT 0.407 0.700 0.480 0.761 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.149 0.706 1.168 0.761 ;
      RECT 1.149 0.520 1.164 0.601 ;
      RECT 1.088 0.520 1.149 0.761 ;
      RECT 1.074 0.520 1.088 0.601 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.864 0.505 1.013 0.633 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.782 0.706 0.818 0.761 ;
      RECT 0.721 0.536 0.782 0.761 ;
      RECT 0.672 0.536 0.721 0.617 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.520 -0.080 1.400 0.080 ;
      RECT 0.430 -0.080 0.520 0.289 ;
      RECT 0.138 -0.080 0.430 0.080 ;
      RECT 0.048 -0.080 0.138 0.330 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.217 1.120 1.400 1.280 ;
      RECT 1.127 1.078 1.217 1.280 ;
      RECT 0.138 1.120 1.127 1.280 ;
      RECT 0.048 0.800 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.002 0.201 1.092 0.304 ;
      RECT 0.711 0.201 1.002 0.256 ;
      RECT 0.681 0.201 0.711 0.350 ;
      RECT 0.650 0.201 0.681 0.413 ;
      RECT 0.620 0.269 0.650 0.413 ;
      RECT 0.329 0.358 0.620 0.413 ;
      RECT 0.268 0.263 0.329 0.413 ;
      RECT 0.239 0.263 0.268 0.344 ;
  END
END OAI33X1

MACRO OAI32X4
  CLASS CORE ;
  FOREIGN OAI32X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.361 0.433 1.402 0.767 ;
      RECT 1.298 0.348 1.361 0.767 ;
      RECT 1.211 0.348 1.298 0.402 ;
      RECT 1.139 0.688 1.298 0.743 ;
      RECT 1.118 0.321 1.211 0.402 ;
      RECT 1.043 0.688 1.139 0.769 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.567 0.142 0.740 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.955 0.391 1.049 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.884 0.567 1.042 0.633 ;
      RECT 0.791 0.526 0.884 0.633 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.695 0.706 0.841 0.761 ;
      RECT 0.633 0.527 0.695 0.761 ;
      RECT 0.603 0.527 0.633 0.608 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.385 0.567 0.502 0.717 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.396 -0.080 1.800 0.080 ;
      RECT 1.304 -0.080 1.396 0.122 ;
      RECT 1.006 -0.080 1.304 0.080 ;
      RECT 0.914 -0.080 1.006 0.122 ;
      RECT 0.698 -0.080 0.914 0.080 ;
      RECT 0.605 -0.080 0.698 0.122 ;
      RECT 0.000 -0.080 0.605 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.358 1.120 1.800 1.280 ;
      RECT 1.265 0.989 1.358 1.280 ;
      RECT 0.961 1.120 1.265 1.280 ;
      RECT 0.869 0.989 0.961 1.280 ;
      RECT 0.142 1.120 0.869 1.280 ;
      RECT 0.049 1.078 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.591 0.194 1.654 0.812 ;
      RECT 1.512 0.194 1.591 0.304 ;
      RECT 1.465 0.605 1.527 0.880 ;
      RECT 1.039 0.194 1.512 0.249 ;
      RECT 0.447 0.825 1.465 0.880 ;
      RECT 1.105 0.457 1.197 0.538 ;
      RECT 1.039 0.457 1.105 0.512 ;
      RECT 0.976 0.194 1.039 0.512 ;
      RECT 0.758 0.300 0.851 0.381 ;
      RECT 0.491 0.313 0.758 0.368 ;
      RECT 0.398 0.300 0.491 0.381 ;
      RECT 0.355 0.808 0.447 0.889 ;
      RECT 0.267 0.808 0.355 0.863 ;
      RECT 0.267 0.300 0.295 0.381 ;
      RECT 0.205 0.300 0.267 0.863 ;
      RECT 0.202 0.300 0.205 0.381 ;
  END
END OAI32X4

MACRO OAI32X1
  CLASS CORE ;
  FOREIGN OAI32X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.360 1.240 0.876 ;
      RECT 1.154 0.360 1.175 0.439 ;
      RECT 0.568 0.821 1.175 0.876 ;
      RECT 0.957 0.360 1.154 0.414 ;
      RECT 0.861 0.314 0.957 0.414 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.929 0.487 1.075 0.640 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.706 0.868 0.761 ;
      RECT 0.734 0.542 0.799 0.761 ;
      RECT 0.703 0.542 0.734 0.623 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.567 0.149 0.711 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.332 0.456 0.402 0.511 ;
      RECT 0.246 0.456 0.332 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.432 0.613 0.560 0.761 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.552 -0.080 1.300 0.080 ;
      RECT 0.456 -0.080 0.552 0.277 ;
      RECT 0.146 -0.080 0.456 0.080 ;
      RECT 0.051 -0.080 0.146 0.290 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.035 1.120 1.300 1.280 ;
      RECT 0.940 1.065 1.035 1.280 ;
      RECT 0.146 1.120 0.940 1.280 ;
      RECT 0.051 1.002 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.064 0.205 1.159 0.305 ;
      RECT 0.754 0.205 1.064 0.260 ;
      RECT 0.723 0.205 0.754 0.345 ;
      RECT 0.689 0.205 0.723 0.401 ;
      RECT 0.658 0.264 0.689 0.401 ;
      RECT 0.349 0.346 0.658 0.401 ;
      RECT 0.284 0.257 0.349 0.401 ;
      RECT 0.253 0.257 0.284 0.338 ;
  END
END OAI32X1

MACRO OAI31X1
  CLASS CORE ;
  FOREIGN OAI31X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.976 0.236 1.040 0.845 ;
      RECT 0.956 0.236 0.976 0.306 ;
      RECT 0.956 0.761 0.976 0.845 ;
      RECT 0.872 0.236 0.956 0.290 ;
      RECT 0.572 0.790 0.956 0.845 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.793 0.440 0.885 0.627 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.481 0.144 0.633 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.433 0.411 0.507 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.486 0.549 0.603 0.651 ;
      RECT 0.426 0.570 0.486 0.627 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.567 -0.080 1.100 0.080 ;
      RECT 0.556 -0.080 0.567 0.087 ;
      RECT 0.461 -0.080 0.556 0.122 ;
      RECT 0.450 -0.080 0.461 0.087 ;
      RECT 0.144 -0.080 0.450 0.080 ;
      RECT 0.050 -0.080 0.144 0.275 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.822 1.120 1.100 1.280 ;
      RECT 0.728 1.078 0.822 1.280 ;
      RECT 0.144 1.120 0.728 1.280 ;
      RECT 0.050 0.925 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.250 0.296 0.767 0.351 ;
  END
END OAI31X1

MACRO OAI2BB2X4
  CLASS CORE ;
  FOREIGN OAI2BB2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.524 0.279 2.553 0.360 ;
      RECT 2.463 0.192 2.524 0.492 ;
      RECT 1.480 0.192 2.463 0.246 ;
      RECT 2.390 0.437 2.463 0.492 ;
      RECT 2.290 0.433 2.390 0.826 ;
      RECT 1.620 0.745 2.290 0.826 ;
      RECT 1.559 0.701 1.620 0.826 ;
      RECT 1.175 0.701 1.559 0.756 ;
      RECT 1.391 0.157 1.480 0.246 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.850 0.565 1.908 0.620 ;
      RECT 1.831 0.565 1.850 0.629 ;
      RECT 1.790 0.565 1.831 0.646 ;
      RECT 1.770 0.574 1.790 0.646 ;
      RECT 0.997 0.592 1.770 0.646 ;
      RECT 0.907 0.533 0.997 0.646 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.197 0.456 2.230 0.573 ;
      RECT 2.136 0.456 2.197 0.627 ;
      RECT 1.710 0.456 2.136 0.511 ;
      RECT 1.694 0.456 1.710 0.530 ;
      RECT 1.648 0.456 1.694 0.537 ;
      RECT 1.619 0.475 1.648 0.537 ;
      RECT 1.112 0.482 1.619 0.537 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.339 0.555 0.428 0.636 ;
      RECT 0.289 0.555 0.339 0.633 ;
      RECT 0.217 0.567 0.289 0.633 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.671 0.444 0.746 0.525 ;
      RECT 0.657 0.185 0.671 0.525 ;
      RECT 0.611 0.185 0.657 0.499 ;
      RECT 0.303 0.185 0.611 0.239 ;
      RECT 0.243 0.185 0.303 0.481 ;
      RECT 0.230 0.426 0.243 0.481 ;
      RECT 0.160 0.426 0.230 0.500 ;
      RECT 0.071 0.426 0.160 0.507 ;
      RECT 0.056 0.439 0.071 0.494 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.185 -0.080 2.600 0.080 ;
      RECT 2.096 -0.080 2.185 0.122 ;
      RECT 1.827 -0.080 2.096 0.080 ;
      RECT 1.737 -0.080 1.827 0.122 ;
      RECT 1.112 -0.080 1.737 0.080 ;
      RECT 0.731 -0.080 1.112 0.122 ;
      RECT 0.137 -0.080 0.731 0.080 ;
      RECT 0.047 -0.080 0.137 0.275 ;
      RECT 0.000 -0.080 0.047 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.542 1.120 2.600 1.280 ;
      RECT 2.453 1.078 2.542 1.280 ;
      RECT 1.995 1.120 2.453 1.280 ;
      RECT 1.905 1.078 1.995 1.280 ;
      RECT 1.448 1.120 1.905 1.280 ;
      RECT 1.359 1.078 1.448 1.280 ;
      RECT 0.918 1.120 1.359 1.280 ;
      RECT 0.829 1.078 0.918 1.280 ;
      RECT 0.523 1.120 0.829 1.280 ;
      RECT 0.433 1.078 0.523 1.280 ;
      RECT 0.137 1.120 0.433 1.280 ;
      RECT 0.047 0.791 0.137 1.280 ;
      RECT 0.000 1.120 0.047 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.450 0.546 2.540 1.006 ;
      RECT 1.481 0.925 2.450 1.006 ;
      RECT 2.194 0.324 2.364 0.379 ;
      RECT 2.134 0.324 2.194 0.401 ;
      RECT 1.312 0.346 2.134 0.401 ;
      RECT 1.392 0.814 1.481 1.006 ;
      RECT 1.110 0.814 1.392 0.895 ;
      RECT 1.223 0.331 1.312 0.412 ;
      RECT 0.961 0.346 1.223 0.401 ;
      RECT 1.020 0.736 1.110 0.895 ;
      RECT 0.549 0.736 1.020 0.817 ;
      RECT 0.872 0.331 0.961 0.412 ;
      RECT 0.488 0.320 0.549 0.817 ;
      RECT 0.473 0.320 0.488 0.375 ;
      RECT 0.236 0.736 0.488 0.817 ;
      RECT 0.383 0.294 0.473 0.375 ;
  END
END OAI2BB2X4

MACRO OAI2BB2X2
  CLASS CORE ;
  FOREIGN OAI2BB2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.679 0.406 1.741 0.923 ;
      RECT 1.231 0.406 1.679 0.461 ;
      RECT 1.316 0.868 1.679 0.923 ;
      RECT 1.223 0.868 1.316 0.949 ;
      RECT 1.169 0.301 1.231 0.461 ;
      RECT 0.901 0.868 1.223 0.923 ;
      RECT 1.102 0.301 1.169 0.356 ;
      RECT 0.809 0.868 0.901 0.949 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 0.626 1.583 0.761 ;
      RECT 1.520 0.626 1.541 0.801 ;
      RECT 1.478 0.706 1.520 0.801 ;
      RECT 1.240 0.746 1.478 0.801 ;
      RECT 1.177 0.632 1.240 0.801 ;
      RECT 1.118 0.632 1.177 0.706 ;
      RECT 0.649 0.632 1.118 0.687 ;
      RECT 0.586 0.529 0.649 0.687 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.370 0.637 1.415 0.692 ;
      RECT 1.308 0.520 1.370 0.692 ;
      RECT 0.920 0.520 1.308 0.575 ;
      RECT 0.858 0.439 0.920 0.575 ;
      RECT 0.779 0.439 0.858 0.494 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.567 0.398 0.690 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.388 0.207 0.512 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.544 -0.080 1.800 0.080 ;
      RECT 1.451 -0.080 1.544 0.122 ;
      RECT 0.791 -0.080 1.451 0.080 ;
      RECT 0.698 -0.080 0.791 0.122 ;
      RECT 0.142 -0.080 0.698 0.080 ;
      RECT 0.049 -0.080 0.142 0.289 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.676 1.120 1.800 1.280 ;
      RECT 1.583 1.078 1.676 1.280 ;
      RECT 1.109 1.120 1.583 1.280 ;
      RECT 1.016 1.078 1.109 1.280 ;
      RECT 0.552 1.120 1.016 1.280 ;
      RECT 0.460 0.902 0.552 1.280 ;
      RECT 0.160 1.120 0.460 1.280 ;
      RECT 0.067 0.832 0.160 1.280 ;
      RECT 0.000 1.120 0.067 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.658 0.225 1.751 0.306 ;
      RECT 1.391 0.251 1.658 0.306 ;
      RECT 1.360 0.251 1.391 0.351 ;
      RECT 1.297 0.185 1.360 0.351 ;
      RECT 0.998 0.185 1.297 0.239 ;
      RECT 0.524 0.742 1.004 0.796 ;
      RECT 0.905 0.185 0.998 0.265 ;
      RECT 0.694 0.211 0.905 0.265 ;
      RECT 0.631 0.211 0.694 0.377 ;
      RECT 0.545 0.323 0.631 0.377 ;
      RECT 0.483 0.449 0.524 0.832 ;
      RECT 0.483 0.156 0.502 0.211 ;
      RECT 0.461 0.156 0.483 0.832 ;
      RECT 0.391 0.156 0.461 0.504 ;
      RECT 0.356 0.777 0.461 0.832 ;
      RECT 0.263 0.777 0.356 0.864 ;
  END
END OAI2BB2X2

MACRO OAI2BB2X1
  CLASS CORE ;
  FOREIGN OAI2BB2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.232 0.439 1.240 0.494 ;
      RECT 1.168 0.250 1.232 0.852 ;
      RECT 1.137 0.250 1.168 0.331 ;
      RECT 1.154 0.761 1.168 0.852 ;
      RECT 0.810 0.798 1.154 0.852 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.570 0.514 0.703 0.633 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.768 0.433 0.889 0.595 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.234 0.500 0.342 0.633 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.392 0.169 0.507 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.827 -0.080 1.300 0.080 ;
      RECT 0.732 -0.080 0.827 0.212 ;
      RECT 0.146 -0.080 0.732 0.080 ;
      RECT 0.051 -0.080 0.146 0.122 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.120 1.120 1.300 1.280 ;
      RECT 1.024 1.078 1.120 1.280 ;
      RECT 0.563 1.120 1.024 1.280 ;
      RECT 0.467 1.078 0.563 1.280 ;
      RECT 0.197 1.120 0.467 1.280 ;
      RECT 0.181 1.078 0.197 1.280 ;
      RECT 0.117 1.065 0.181 1.280 ;
      RECT 0.101 1.078 0.117 1.280 ;
      RECT 0.000 1.120 0.101 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.017 0.438 1.082 0.743 ;
      RECT 0.999 0.188 1.030 0.269 ;
      RECT 0.471 0.688 1.017 0.743 ;
      RECT 0.934 0.188 0.999 0.337 ;
      RECT 0.613 0.282 0.934 0.337 ;
      RECT 0.549 0.156 0.613 0.337 ;
      RECT 0.518 0.156 0.549 0.211 ;
      RECT 0.471 0.310 0.473 0.390 ;
      RECT 0.407 0.310 0.471 0.781 ;
      RECT 0.377 0.310 0.407 0.390 ;
      RECT 0.366 0.726 0.407 0.781 ;
      RECT 0.270 0.726 0.366 0.807 ;
  END
END OAI2BB2X1

MACRO OAI2BB1X4
  CLASS CORE ;
  FOREIGN OAI2BB1X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.620 0.170 1.669 0.251 ;
      RECT 1.582 0.170 1.620 0.621 ;
      RECT 1.561 0.170 1.582 0.900 ;
      RECT 1.557 0.183 1.561 0.900 ;
      RECT 1.320 0.183 1.557 0.238 ;
      RECT 1.478 0.567 1.557 0.900 ;
      RECT 1.139 0.701 1.478 0.756 ;
      RECT 1.309 0.170 1.320 0.238 ;
      RECT 1.216 0.170 1.309 0.251 ;
      RECT 1.016 0.688 1.139 0.769 ;
      RECT 0.779 0.701 1.016 0.756 ;
      RECT 0.760 0.701 0.779 0.769 ;
      RECT 0.667 0.688 0.760 0.769 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.578 0.539 0.824 0.633 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.481 0.142 0.633 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.331 0.539 0.502 0.633 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.840 -0.080 1.800 0.080 ;
      RECT 0.747 -0.080 0.840 0.212 ;
      RECT 0.491 -0.080 0.747 0.080 ;
      RECT 0.398 -0.080 0.491 0.212 ;
      RECT 0.000 -0.080 0.398 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.283 1.120 1.800 1.280 ;
      RECT 1.190 0.877 1.283 1.280 ;
      RECT 0.934 1.120 1.190 1.280 ;
      RECT 0.841 0.877 0.934 1.280 ;
      RECT 0.567 1.120 0.841 1.280 ;
      RECT 0.475 0.944 0.567 1.280 ;
      RECT 0.142 1.120 0.475 1.280 ;
      RECT 0.049 0.747 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.402 0.319 1.495 0.424 ;
      RECT 1.065 0.525 1.414 0.606 ;
      RECT 1.047 0.319 1.402 0.374 ;
      RECT 0.972 0.525 1.065 0.580 ;
      RECT 0.955 0.280 1.047 0.374 ;
      RECT 0.910 0.430 0.972 0.580 ;
      RECT 0.650 0.319 0.955 0.374 ;
      RECT 0.267 0.430 0.910 0.485 ;
      RECT 0.588 0.319 0.650 0.375 ;
      RECT 0.573 0.320 0.588 0.375 ;
      RECT 0.267 0.732 0.349 1.037 ;
      RECT 0.256 0.289 0.267 1.037 ;
      RECT 0.205 0.289 0.256 0.788 ;
      RECT 0.142 0.289 0.205 0.344 ;
      RECT 0.049 0.151 0.142 0.344 ;
  END
END OAI2BB1X4

MACRO OAI2BB1X2
  CLASS CORE ;
  FOREIGN OAI2BB1X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.033 0.292 1.054 0.627 ;
      RECT 0.989 0.292 1.033 0.731 ;
      RECT 0.889 0.292 0.989 0.346 ;
      RECT 0.968 0.573 0.989 0.731 ;
      RECT 0.917 0.676 0.968 0.731 ;
      RECT 0.822 0.676 0.917 0.757 ;
      RECT 0.794 0.265 0.889 0.346 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.535 0.379 0.703 0.507 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.060 0.400 0.165 0.533 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.423 0.567 0.568 0.633 ;
      RECT 0.359 0.542 0.423 0.633 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 -0.080 1.300 0.080 ;
      RECT 1.154 -0.080 1.249 0.289 ;
      RECT 0.518 -0.080 1.154 0.080 ;
      RECT 0.422 -0.080 0.518 0.289 ;
      RECT 0.000 -0.080 0.422 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.109 1.120 1.300 1.280 ;
      RECT 1.013 1.078 1.109 1.280 ;
      RECT 0.737 1.120 1.013 1.280 ;
      RECT 0.642 0.972 0.737 1.280 ;
      RECT 0.298 1.120 0.642 1.280 ;
      RECT 0.203 1.078 0.298 1.280 ;
      RECT 0.000 1.120 0.203 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.833 0.468 0.864 0.549 ;
      RECT 0.768 0.468 0.833 0.621 ;
      RECT 0.756 0.567 0.768 0.621 ;
      RECT 0.691 0.567 0.756 0.823 ;
      RECT 0.523 0.768 0.691 0.823 ;
      RECT 0.428 0.768 0.523 0.849 ;
      RECT 0.294 0.768 0.428 0.823 ;
      RECT 0.229 0.280 0.294 0.823 ;
      RECT 0.146 0.280 0.229 0.335 ;
      RECT 0.051 0.254 0.146 0.335 ;
  END
END OAI2BB1X2

MACRO OAI2BB1X1
  CLASS CORE ;
  FOREIGN OAI2BB1X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.798 0.343 0.860 0.913 ;
      RECT 0.758 0.343 0.798 0.424 ;
      RECT 0.779 0.839 0.798 0.913 ;
      RECT 0.678 0.858 0.779 0.913 ;
      RECT 0.585 0.858 0.678 0.939 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.526 0.566 0.640 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.142 0.612 0.185 0.693 ;
      RECT 0.038 0.612 0.142 0.767 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.170 0.424 0.322 0.532 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.513 -0.080 0.900 0.080 ;
      RECT 0.420 -0.080 0.513 0.122 ;
      RECT 0.000 -0.080 0.420 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.830 1.120 0.900 1.280 ;
      RECT 0.815 1.078 0.830 1.280 ;
      RECT 0.753 1.065 0.815 1.280 ;
      RECT 0.738 1.078 0.753 1.280 ;
      RECT 0.469 1.120 0.738 1.280 ;
      RECT 0.049 1.078 0.469 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.695 0.500 0.735 0.583 ;
      RECT 0.633 0.235 0.695 0.804 ;
      RECT 0.142 0.235 0.633 0.289 ;
      RECT 0.305 0.749 0.633 0.804 ;
      RECT 0.213 0.749 0.305 0.843 ;
      RECT 0.049 0.223 0.142 0.304 ;
  END
END OAI2BB1X1

MACRO OAI22X4
  CLASS CORE ;
  FOREIGN OAI22X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.440 0.433 2.462 0.767 ;
      RECT 2.378 0.158 2.440 0.767 ;
      RECT 1.326 0.158 2.378 0.213 ;
      RECT 2.359 0.433 2.378 0.767 ;
      RECT 2.229 0.702 2.359 0.757 ;
      RECT 2.137 0.702 2.229 0.927 ;
      RECT 2.085 0.702 2.137 0.767 ;
      RECT 1.537 0.702 2.085 0.757 ;
      RECT 1.445 0.702 1.537 0.927 ;
      RECT 1.370 0.702 1.445 0.767 ;
      RECT 0.844 0.702 1.370 0.757 ;
      RECT 0.752 0.702 0.844 0.927 ;
      RECT 0.152 0.702 0.752 0.757 ;
      RECT 0.060 0.702 0.152 0.926 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.032 0.537 1.094 0.639 ;
      RECT 0.567 0.585 1.032 0.639 ;
      RECT 0.476 0.550 0.567 0.639 ;
      RECT 0.415 0.550 0.476 0.627 ;
      RECT 0.341 0.550 0.415 0.605 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.760 0.449 0.920 0.530 ;
      RECT 0.687 0.440 0.760 0.530 ;
      RECT 0.120 0.440 0.687 0.495 ;
      RECT 0.058 0.440 0.120 0.627 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.907 0.449 1.937 0.530 ;
      RECT 1.845 0.440 1.907 0.530 ;
      RECT 1.353 0.440 1.845 0.495 ;
      RECT 1.353 0.563 1.370 0.627 ;
      RECT 1.308 0.440 1.353 0.627 ;
      RECT 1.291 0.440 1.308 0.618 ;
      RECT 1.199 0.537 1.291 0.618 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.117 0.537 2.179 0.639 ;
      RECT 2.085 0.567 2.117 0.639 ;
      RECT 1.748 0.585 2.085 0.639 ;
      RECT 1.686 0.550 1.748 0.639 ;
      RECT 1.665 0.550 1.686 0.627 ;
      RECT 1.494 0.550 1.665 0.605 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.028 -0.080 2.500 0.080 ;
      RECT 0.936 -0.080 1.028 0.211 ;
      RECT 0.682 -0.080 0.936 0.080 ;
      RECT 0.590 -0.080 0.682 0.211 ;
      RECT 0.335 -0.080 0.590 0.080 ;
      RECT 0.244 -0.080 0.335 0.211 ;
      RECT 0.000 -0.080 0.244 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.883 1.120 2.500 1.280 ;
      RECT 1.791 0.932 1.883 1.280 ;
      RECT 1.190 1.120 1.791 1.280 ;
      RECT 1.098 0.932 1.190 1.280 ;
      RECT 0.498 1.120 1.098 1.280 ;
      RECT 0.406 0.932 0.498 1.280 ;
      RECT 0.000 1.120 0.406 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.224 0.269 2.316 0.350 ;
      RECT 2.081 0.295 2.224 0.350 ;
      RECT 2.018 0.295 2.081 0.386 ;
      RECT 1.223 0.331 2.018 0.386 ;
      RECT 1.131 0.217 1.223 0.386 ;
      RECT 0.261 0.331 1.131 0.386 ;
      RECT 0.199 0.330 0.261 0.386 ;
      RECT 0.141 0.330 0.199 0.385 ;
      RECT 0.078 0.217 0.141 0.385 ;
      RECT 0.049 0.217 0.078 0.298 ;
  END
END OAI22X4

MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.976 0.358 1.040 0.894 ;
      RECT 0.956 0.358 0.976 0.439 ;
      RECT 0.511 0.839 0.976 0.894 ;
      RECT 0.767 0.358 0.956 0.413 ;
      RECT 0.703 0.313 0.767 0.413 ;
      RECT 0.672 0.313 0.703 0.394 ;
      RECT 0.417 0.826 0.511 0.907 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.567 0.233 0.655 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.350 0.433 0.444 0.520 ;
      RECT 0.222 0.433 0.350 0.511 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.772 0.585 0.878 0.767 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.575 0.473 0.694 0.633 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.356 -0.080 1.100 0.080 ;
      RECT 0.261 -0.080 0.356 0.122 ;
      RECT 0.000 -0.080 0.261 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.878 1.120 1.100 1.280 ;
      RECT 0.783 1.078 0.878 1.280 ;
      RECT 0.144 1.120 0.783 1.280 ;
      RECT 0.050 1.078 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.936 0.223 0.967 0.304 ;
      RECT 0.872 0.204 0.936 0.304 ;
      RECT 0.567 0.204 0.872 0.258 ;
      RECT 0.503 0.204 0.567 0.379 ;
      RECT 0.472 0.298 0.503 0.379 ;
      RECT 0.144 0.311 0.472 0.365 ;
      RECT 0.050 0.298 0.144 0.379 ;
  END
END OAI22X1

MACRO OAI222XL
  CLASS CORE ;
  FOREIGN OAI222XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.282 0.419 1.343 0.894 ;
      RECT 1.188 0.419 1.282 0.474 ;
      RECT 1.148 0.839 1.282 0.894 ;
      RECT 1.151 0.361 1.188 0.474 ;
      RECT 1.090 0.281 1.151 0.474 ;
      RECT 1.058 0.829 1.148 0.910 ;
      RECT 1.061 0.281 1.090 0.362 ;
      RECT 0.993 0.833 1.058 0.900 ;
      RECT 0.435 0.842 0.993 0.896 ;
      RECT 0.345 0.829 0.435 0.910 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.860 0.507 1.013 0.633 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.086 0.615 1.214 0.767 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.567 0.138 0.715 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.413 0.337 0.558 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.562 0.577 0.676 0.768 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.353 0.639 0.488 0.767 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 -0.080 1.400 0.080 ;
      RECT 0.345 -0.080 0.435 0.122 ;
      RECT 0.138 -0.080 0.345 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.791 1.120 1.400 1.280 ;
      RECT 0.701 1.078 0.791 1.280 ;
      RECT 0.138 1.120 0.701 1.280 ;
      RECT 0.048 1.078 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.313 0.281 1.342 0.362 ;
      RECT 1.252 0.155 1.313 0.362 ;
      RECT 0.960 0.155 1.252 0.210 ;
      RECT 0.899 0.155 0.960 0.362 ;
      RECT 0.870 0.281 0.899 0.362 ;
      RECT 0.679 0.252 0.769 0.362 ;
      RECT 0.286 0.252 0.679 0.307 ;
      RECT 0.196 0.252 0.286 0.333 ;
  END
END OAI222XL

MACRO OAI221XL
  CLASS CORE ;
  FOREIGN OAI221XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.258 1.240 0.920 ;
      RECT 1.095 0.258 1.175 0.339 ;
      RECT 0.990 0.865 1.175 0.920 ;
      RECT 0.895 0.865 0.990 0.946 ;
      RECT 0.461 0.865 0.895 0.920 ;
      RECT 0.366 0.865 0.461 0.946 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.968 0.521 1.075 0.654 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.640 0.146 0.821 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.187 0.433 0.359 0.550 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.803 0.700 0.868 0.761 ;
      RECT 0.718 0.700 0.803 0.755 ;
      RECT 0.622 0.639 0.718 0.755 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.516 0.642 0.519 0.779 ;
      RECT 0.421 0.640 0.516 0.779 ;
      RECT 0.336 0.642 0.421 0.779 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.461 -0.080 1.300 0.080 ;
      RECT 0.366 -0.080 0.461 0.122 ;
      RECT 0.146 -0.080 0.366 0.080 ;
      RECT 0.051 -0.080 0.146 0.122 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.777 1.120 1.300 1.280 ;
      RECT 0.681 1.078 0.777 1.280 ;
      RECT 0.146 1.120 0.681 1.280 ;
      RECT 0.051 1.078 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.786 0.339 0.817 0.420 ;
      RECT 0.722 0.252 0.786 0.420 ;
      RECT 0.304 0.252 0.722 0.307 ;
      RECT 0.208 0.252 0.304 0.333 ;
  END
END OAI221XL

MACRO OAI221X4
  CLASS CORE ;
  FOREIGN OAI221X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.740 0.433 1.780 0.767 ;
      RECT 1.708 0.290 1.740 0.767 ;
      RECT 1.682 0.154 1.708 0.767 ;
      RECT 1.676 0.154 1.682 0.975 ;
      RECT 1.614 0.154 1.676 0.346 ;
      RECT 1.675 0.433 1.676 0.975 ;
      RECT 1.588 0.670 1.675 0.975 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.948 0.560 1.052 0.696 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.654 0.165 0.790 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.220 0.407 0.405 0.517 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.787 0.573 0.850 0.633 ;
      RECT 0.704 0.579 0.787 0.633 ;
      RECT 0.640 0.579 0.704 0.735 ;
      RECT 0.610 0.654 0.640 0.735 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.402 0.651 0.518 0.789 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.906 -0.080 2.000 0.080 ;
      RECT 1.813 -0.080 1.906 0.323 ;
      RECT 1.510 -0.080 1.813 0.080 ;
      RECT 1.416 -0.080 1.510 0.324 ;
      RECT 0.452 -0.080 1.416 0.080 ;
      RECT 0.358 -0.080 0.452 0.122 ;
      RECT 0.143 -0.080 0.358 0.080 ;
      RECT 0.050 -0.080 0.143 0.122 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.880 1.120 2.000 1.280 ;
      RECT 1.787 0.876 1.880 1.280 ;
      RECT 1.472 1.120 1.787 1.280 ;
      RECT 1.379 1.078 1.472 1.280 ;
      RECT 1.164 1.120 1.379 1.280 ;
      RECT 1.070 1.078 1.164 1.280 ;
      RECT 0.760 1.120 1.070 1.280 ;
      RECT 0.667 1.078 0.760 1.280 ;
      RECT 0.143 1.120 0.667 1.280 ;
      RECT 0.050 1.078 0.143 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.475 0.457 1.569 0.538 ;
      RECT 1.379 0.470 1.475 0.538 ;
      RECT 1.318 0.402 1.379 0.933 ;
      RECT 1.315 0.402 1.318 0.946 ;
      RECT 1.311 0.402 1.315 0.457 ;
      RECT 1.225 0.865 1.315 0.946 ;
      RECT 1.248 0.215 1.311 0.457 ;
      RECT 1.179 0.544 1.252 0.625 ;
      RECT 1.218 0.215 1.248 0.296 ;
      RECT 1.116 0.385 1.179 0.810 ;
      RECT 1.069 0.385 1.116 0.465 ;
      RECT 0.971 0.755 1.116 0.810 ;
      RECT 0.908 0.755 0.971 0.944 ;
      RECT 0.358 0.863 0.908 0.944 ;
      RECT 0.705 0.298 0.799 0.419 ;
      RECT 0.298 0.298 0.705 0.352 ;
      RECT 0.204 0.271 0.298 0.352 ;
  END
END OAI221X4

MACRO OAI221X2
  CLASS CORE ;
  FOREIGN OAI221X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.976 0.345 2.032 0.830 ;
      RECT 1.970 0.318 1.976 0.830 ;
      RECT 1.914 0.318 1.970 0.440 ;
      RECT 1.732 0.775 1.970 0.830 ;
      RECT 1.716 0.775 1.732 0.839 ;
      RECT 1.654 0.775 1.716 0.904 ;
      RECT 1.624 0.823 1.654 0.904 ;
      RECT 1.169 0.839 1.624 0.894 ;
      RECT 1.078 0.839 1.169 0.920 ;
      RECT 1.003 0.839 1.078 0.900 ;
      RECT 0.483 0.839 1.003 0.894 ;
      RECT 0.391 0.839 0.483 0.920 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.647 0.567 1.903 0.633 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.204 0.552 0.740 0.607 ;
      RECT 0.113 0.546 0.204 0.627 ;
      RECT 0.058 0.573 0.113 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.473 0.662 0.547 0.743 ;
      RECT 0.411 0.662 0.473 0.761 ;
      RECT 0.327 0.662 0.411 0.743 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.319 0.562 1.512 0.617 ;
      RECT 1.257 0.552 1.319 0.617 ;
      RECT 1.004 0.552 1.257 0.607 ;
      RECT 0.954 0.552 1.004 0.627 ;
      RECT 0.942 0.552 0.954 0.640 ;
      RECT 0.863 0.560 0.942 0.640 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.196 0.700 1.240 0.767 ;
      RECT 1.104 0.662 1.196 0.767 ;
      RECT 1.024 0.700 1.104 0.767 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.869 -0.080 2.300 0.080 ;
      RECT 0.777 -0.080 0.869 0.211 ;
      RECT 0.483 -0.080 0.777 0.080 ;
      RECT 0.391 -0.080 0.483 0.211 ;
      RECT 0.139 -0.080 0.391 0.080 ;
      RECT 0.048 -0.080 0.139 0.211 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.909 1.120 2.300 1.280 ;
      RECT 1.817 0.900 1.909 1.280 ;
      RECT 1.512 1.120 1.817 1.280 ;
      RECT 1.421 0.984 1.512 1.280 ;
      RECT 0.826 1.120 1.421 1.280 ;
      RECT 0.734 0.984 0.826 1.280 ;
      RECT 0.139 1.120 0.734 1.280 ;
      RECT 0.048 0.929 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.783 0.193 2.162 0.248 ;
      RECT 1.721 0.158 1.783 0.327 ;
      RECT 0.965 0.158 1.721 0.213 ;
      RECT 1.228 0.302 1.604 0.357 ;
      RECT 1.137 0.302 1.228 0.399 ;
      RECT 0.676 0.302 1.137 0.357 ;
      RECT 0.646 0.217 0.676 0.357 ;
      RECT 0.584 0.217 0.646 0.373 ;
      RECT 0.311 0.318 0.584 0.373 ;
      RECT 0.220 0.318 0.311 0.399 ;
  END
END OAI221X2

MACRO OAI221X1
  CLASS CORE ;
  FOREIGN OAI221X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.310 0.829 1.358 0.910 ;
      RECT 1.249 0.282 1.310 0.910 ;
      RECT 1.204 0.282 1.249 0.363 ;
      RECT 0.398 0.829 1.249 0.910 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.017 0.533 1.188 0.640 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.567 0.223 0.655 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.399 0.412 0.500 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.673 0.567 0.838 0.671 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.375 0.560 0.581 0.673 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.541 -0.080 1.400 0.080 ;
      RECT 0.451 -0.080 0.541 0.122 ;
      RECT 0.138 -0.080 0.451 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.838 1.120 1.400 1.280 ;
      RECT 0.823 1.078 0.838 1.280 ;
      RECT 0.762 1.065 0.823 1.280 ;
      RECT 0.748 1.078 0.762 1.280 ;
      RECT 0.138 1.120 0.748 1.280 ;
      RECT 0.048 1.078 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.013 0.337 1.103 0.418 ;
      RECT 0.721 0.363 1.013 0.418 ;
      RECT 0.822 0.226 0.912 0.307 ;
      RECT 0.339 0.226 0.822 0.281 ;
      RECT 0.631 0.345 0.721 0.426 ;
      RECT 0.249 0.226 0.339 0.307 ;
  END
END OAI221X1

MACRO OAI21XL
  CLASS CORE ;
  FOREIGN OAI21XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.643 0.439 0.650 0.915 ;
      RECT 0.589 0.161 0.643 0.915 ;
      RECT 0.582 0.161 0.589 0.494 ;
      RECT 0.477 0.861 0.589 0.915 ;
      RECT 0.546 0.161 0.582 0.215 ;
      RECT 0.387 0.848 0.477 0.929 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.640 0.528 0.767 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.048 0.433 0.138 0.618 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.293 0.479 0.388 0.571 ;
      RECT 0.232 0.439 0.293 0.571 ;
      RECT 0.212 0.479 0.232 0.571 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.286 -0.080 0.700 0.080 ;
      RECT 0.196 -0.080 0.286 0.122 ;
      RECT 0.000 -0.080 0.196 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.626 1.120 0.700 1.280 ;
      RECT 0.536 1.078 0.626 1.280 ;
      RECT 0.138 1.120 0.536 1.280 ;
      RECT 0.048 0.910 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.459 0.332 0.488 0.413 ;
      RECT 0.398 0.296 0.459 0.413 ;
      RECT 0.138 0.296 0.398 0.351 ;
      RECT 0.048 0.296 0.138 0.377 ;
  END
END OAI21XL

MACRO OAI21X4
  CLASS CORE ;
  FOREIGN OAI21X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.780 0.313 1.809 0.440 ;
      RECT 1.715 0.313 1.780 0.767 ;
      RECT 1.675 0.331 1.715 0.767 ;
      RECT 1.329 0.331 1.675 0.386 ;
      RECT 1.576 0.708 1.675 0.763 ;
      RECT 1.482 0.695 1.576 0.776 ;
      RECT 1.223 0.708 1.482 0.763 ;
      RECT 1.193 0.695 1.223 0.776 ;
      RECT 1.129 0.695 1.193 0.865 ;
      RECT 0.496 0.811 1.129 0.865 ;
      RECT 0.402 0.798 0.496 0.879 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.262 0.560 1.488 0.640 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.788 0.550 0.937 0.605 ;
      RECT 0.752 0.550 0.788 0.633 ;
      RECT 0.689 0.550 0.752 0.743 ;
      RECT 0.209 0.688 0.689 0.743 ;
      RECT 0.146 0.533 0.209 0.743 ;
      RECT 0.131 0.533 0.146 0.633 ;
      RECT 0.116 0.533 0.131 0.627 ;
      RECT 0.059 0.573 0.116 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.091 0.505 1.121 0.586 ;
      RECT 1.028 0.440 1.091 0.586 ;
      RECT 0.584 0.440 1.028 0.495 ;
      RECT 0.521 0.440 0.584 0.614 ;
      RECT 0.492 0.533 0.521 0.614 ;
      RECT 0.423 0.533 0.492 0.627 ;
      RECT 0.336 0.533 0.423 0.614 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.047 -0.080 2.000 0.080 ;
      RECT 0.953 -0.080 1.047 0.211 ;
      RECT 0.694 -0.080 0.953 0.080 ;
      RECT 0.601 -0.080 0.694 0.211 ;
      RECT 0.342 -0.080 0.601 0.080 ;
      RECT 0.248 -0.080 0.342 0.211 ;
      RECT 0.000 -0.080 0.248 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.753 1.120 2.000 1.280 ;
      RECT 1.660 0.883 1.753 1.280 ;
      RECT 1.399 1.120 1.660 1.280 ;
      RECT 1.306 0.883 1.399 1.280 ;
      RECT 0.860 1.120 1.306 1.280 ;
      RECT 0.766 0.947 0.860 1.280 ;
      RECT 0.143 1.120 0.766 1.280 ;
      RECT 0.050 0.847 0.143 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.506 0.150 1.599 0.231 ;
      RECT 1.247 0.163 1.506 0.218 ;
      RECT 1.216 0.150 1.247 0.231 ;
      RECT 1.153 0.150 1.216 0.386 ;
      RECT 0.143 0.331 1.153 0.386 ;
      RECT 0.080 0.226 0.143 0.386 ;
      RECT 0.050 0.226 0.080 0.307 ;
  END
END OAI21X4

MACRO OAI21X2
  CLASS CORE ;
  FOREIGN OAI21X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.283 0.311 1.343 0.920 ;
      RECT 1.282 0.311 1.283 0.946 ;
      RECT 1.114 0.311 1.282 0.365 ;
      RECT 1.151 0.865 1.282 0.946 ;
      RECT 0.838 0.865 1.151 0.920 ;
      RECT 1.053 0.263 1.114 0.365 ;
      RECT 1.023 0.263 1.053 0.344 ;
      RECT 0.748 0.865 0.838 0.946 ;
      RECT 0.138 0.865 0.748 0.920 ;
      RECT 0.048 0.865 0.138 0.946 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 0.551 1.179 0.632 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.614 0.562 0.695 ;
      RECT 0.473 0.614 0.488 0.707 ;
      RECT 0.407 0.614 0.473 0.761 ;
      RECT 0.323 0.614 0.407 0.707 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.711 0.605 0.740 0.686 ;
      RECT 0.650 0.460 0.711 0.686 ;
      RECT 0.232 0.460 0.650 0.514 ;
      RECT 0.119 0.433 0.232 0.514 ;
      RECT 0.118 0.439 0.119 0.514 ;
      RECT 0.057 0.439 0.118 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.732 -0.080 1.400 0.080 ;
      RECT 0.642 -0.080 0.732 0.280 ;
      RECT 0.339 -0.080 0.642 0.080 ;
      RECT 0.249 -0.080 0.339 0.122 ;
      RECT 0.000 -0.080 0.249 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.039 1.120 1.400 1.280 ;
      RECT 0.949 1.078 1.039 1.280 ;
      RECT 0.488 1.120 0.949 1.280 ;
      RECT 0.398 1.078 0.488 1.280 ;
      RECT 0.000 1.120 0.398 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.275 0.175 1.305 0.256 ;
      RECT 1.214 0.154 1.275 0.256 ;
      RECT 0.923 0.154 1.214 0.208 ;
      RECT 0.894 0.154 0.923 0.283 ;
      RECT 0.862 0.154 0.894 0.405 ;
      RECT 0.833 0.202 0.862 0.405 ;
      RECT 0.541 0.350 0.833 0.405 ;
      RECT 0.526 0.223 0.541 0.405 ;
      RECT 0.480 0.221 0.526 0.405 ;
      RECT 0.451 0.221 0.480 0.304 ;
      RECT 0.138 0.221 0.451 0.276 ;
      RECT 0.048 0.195 0.138 0.276 ;
  END
END OAI21X2

MACRO OAI21X1
  CLASS CORE ;
  FOREIGN OAI21X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.780 0.294 0.841 0.915 ;
      RECT 0.779 0.268 0.780 0.915 ;
      RECT 0.660 0.268 0.779 0.349 ;
      RECT 0.513 0.861 0.779 0.915 ;
      RECT 0.420 0.848 0.513 0.929 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.554 0.560 0.682 0.704 ;
      RECT 0.551 0.560 0.554 0.640 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.164 0.433 0.240 0.500 ;
      RECT 0.071 0.426 0.164 0.507 ;
      RECT 0.038 0.433 0.071 0.500 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.567 0.425 0.633 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.349 -0.080 0.900 0.080 ;
      RECT 0.256 -0.080 0.349 0.122 ;
      RECT 0.000 -0.080 0.256 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.720 1.120 0.900 1.280 ;
      RECT 0.627 1.078 0.720 1.280 ;
      RECT 0.142 1.120 0.627 1.280 ;
      RECT 0.049 0.905 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.541 0.223 0.556 0.304 ;
      RECT 0.464 0.218 0.541 0.304 ;
      RECT 0.142 0.218 0.464 0.273 ;
      RECT 0.049 0.205 0.142 0.286 ;
  END
END OAI21X1

MACRO OAI211X4
  CLASS CORE ;
  FOREIGN OAI211X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.552 0.300 1.562 0.633 ;
      RECT 1.460 0.300 1.552 0.757 ;
      RECT 1.288 0.318 1.460 0.399 ;
      RECT 1.201 0.676 1.460 0.757 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.369 0.426 0.560 0.507 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.673 0.537 0.851 0.662 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.337 0.569 0.366 0.650 ;
      RECT 0.275 0.569 0.337 0.761 ;
      RECT 0.236 0.706 0.275 0.761 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.511 0.186 0.635 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.552 -0.080 1.600 0.080 ;
      RECT 1.460 -0.080 1.552 0.211 ;
      RECT 1.207 -0.080 1.460 0.080 ;
      RECT 1.115 -0.080 1.207 0.211 ;
      RECT 0.318 -0.080 1.115 0.080 ;
      RECT 0.226 -0.080 0.318 0.122 ;
      RECT 0.000 -0.080 0.226 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.465 1.120 1.600 1.280 ;
      RECT 1.374 0.972 1.465 1.280 ;
      RECT 1.121 1.120 1.374 1.280 ;
      RECT 1.029 0.972 1.121 1.280 ;
      RECT 0.700 1.120 1.029 1.280 ;
      RECT 0.404 1.078 0.700 1.280 ;
      RECT 0.000 1.120 0.404 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.139 0.462 1.341 0.543 ;
      RECT 1.077 0.281 1.139 0.902 ;
      RECT 1.002 0.281 1.077 0.336 ;
      RECT 0.916 0.848 1.077 0.902 ;
      RECT 0.986 0.483 1.015 0.564 ;
      RECT 0.940 0.150 1.002 0.336 ;
      RECT 0.924 0.394 0.986 0.793 ;
      RECT 0.910 0.150 0.940 0.231 ;
      RECT 0.851 0.394 0.924 0.449 ;
      RECT 0.646 0.738 0.924 0.793 ;
      RECT 0.824 0.848 0.916 0.929 ;
      RECT 0.789 0.317 0.851 0.449 ;
      RECT 0.760 0.317 0.789 0.398 ;
      RECT 0.617 0.738 0.646 0.819 ;
      RECT 0.555 0.738 0.617 0.933 ;
      RECT 0.140 0.879 0.555 0.933 ;
      RECT 0.404 0.269 0.496 0.350 ;
      RECT 0.140 0.277 0.404 0.332 ;
      RECT 0.048 0.257 0.140 0.338 ;
      RECT 0.048 0.879 0.140 0.960 ;
  END
END OAI211X4

MACRO OAI211X2
  CLASS CORE ;
  FOREIGN OAI211X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.631 0.310 1.694 0.755 ;
      RECT 1.319 0.310 1.631 0.364 ;
      RECT 1.561 0.700 1.631 0.755 ;
      RECT 1.541 0.700 1.561 0.761 ;
      RECT 1.499 0.700 1.541 0.920 ;
      RECT 1.478 0.706 1.499 0.920 ;
      RECT 1.320 0.865 1.478 0.920 ;
      RECT 1.184 0.865 1.320 0.946 ;
      RECT 1.298 0.306 1.319 0.364 ;
      RECT 1.205 0.283 1.298 0.364 ;
      RECT 0.862 0.865 1.184 0.920 ;
      RECT 0.769 0.865 0.862 0.952 ;
      RECT 0.142 0.865 0.769 0.920 ;
      RECT 0.049 0.865 0.142 0.946 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.538 0.419 1.568 0.500 ;
      RECT 1.475 0.419 1.538 0.627 ;
      RECT 1.013 0.573 1.475 0.627 ;
      RECT 0.950 0.460 1.013 0.627 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.364 0.439 1.381 0.494 ;
      RECT 1.140 0.426 1.364 0.507 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.502 0.614 0.578 0.695 ;
      RECT 0.487 0.614 0.502 0.707 ;
      RECT 0.419 0.614 0.487 0.761 ;
      RECT 0.333 0.614 0.419 0.707 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.731 0.605 0.761 0.686 ;
      RECT 0.668 0.460 0.731 0.686 ;
      RECT 0.239 0.460 0.668 0.514 ;
      RECT 0.215 0.433 0.239 0.514 ;
      RECT 0.123 0.426 0.215 0.514 ;
      RECT 0.121 0.439 0.123 0.514 ;
      RECT 0.059 0.439 0.121 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.753 -0.080 1.800 0.080 ;
      RECT 0.660 -0.080 0.753 0.280 ;
      RECT 0.349 -0.080 0.660 0.080 ;
      RECT 0.256 -0.080 0.349 0.122 ;
      RECT 0.000 -0.080 0.256 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.069 1.120 1.800 1.280 ;
      RECT 0.976 1.078 1.069 1.280 ;
      RECT 0.502 1.120 0.976 1.280 ;
      RECT 0.409 1.078 0.502 1.280 ;
      RECT 0.000 1.120 0.409 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.555 0.171 1.647 0.252 ;
      RECT 0.949 0.174 1.555 0.229 ;
      RECT 0.919 0.174 0.949 0.283 ;
      RECT 0.886 0.174 0.919 0.405 ;
      RECT 0.856 0.202 0.886 0.405 ;
      RECT 0.556 0.350 0.856 0.405 ;
      RECT 0.541 0.223 0.556 0.405 ;
      RECT 0.494 0.221 0.541 0.405 ;
      RECT 0.464 0.221 0.494 0.304 ;
      RECT 0.142 0.221 0.464 0.276 ;
      RECT 0.049 0.195 0.142 0.276 ;
  END
END OAI211X2

MACRO OAI211X1
  CLASS CORE ;
  FOREIGN OAI211X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.978 0.298 1.040 0.902 ;
      RECT 0.976 0.271 0.978 0.929 ;
      RECT 0.839 0.271 0.976 0.352 ;
      RECT 0.850 0.848 0.976 0.929 ;
      RECT 0.522 0.848 0.850 0.902 ;
      RECT 0.428 0.848 0.522 0.929 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.564 0.560 0.694 0.704 ;
      RECT 0.561 0.560 0.564 0.640 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.772 0.433 0.878 0.602 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.167 0.433 0.244 0.500 ;
      RECT 0.072 0.426 0.167 0.507 ;
      RECT 0.039 0.433 0.072 0.500 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.567 0.433 0.633 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.356 -0.080 1.100 0.080 ;
      RECT 0.261 -0.080 0.356 0.122 ;
      RECT 0.000 -0.080 0.261 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.733 1.120 1.100 1.280 ;
      RECT 0.639 1.078 0.733 1.280 ;
      RECT 0.144 1.120 0.639 1.280 ;
      RECT 0.050 0.905 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.472 0.205 0.567 0.286 ;
      RECT 0.144 0.218 0.472 0.273 ;
      RECT 0.050 0.205 0.144 0.286 ;
  END
END OAI211X1

MACRO NOR4BBX1
  CLASS CORE ;
  FOREIGN NOR4BBX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.307 0.192 1.368 0.894 ;
      RECT 0.888 0.192 1.307 0.246 ;
      RECT 1.014 0.839 1.307 0.894 ;
      RECT 0.924 0.839 1.014 0.920 ;
      RECT 0.813 0.192 0.888 0.339 ;
      RECT 0.798 0.223 0.813 0.339 ;
      RECT 0.418 0.223 0.798 0.304 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.403 0.573 0.468 0.627 ;
      RECT 0.342 0.393 0.403 0.627 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.620 0.573 0.643 0.627 ;
      RECT 0.559 0.412 0.620 0.627 ;
      RECT 0.505 0.412 0.559 0.493 ;
     END
  END C

  PIN BN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.083 0.542 1.115 0.623 ;
      RECT 1.022 0.542 1.083 0.761 ;
      RECT 0.932 0.700 1.022 0.761 ;
     END
  END BN

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.046 0.438 0.137 0.595 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.090 -0.080 1.400 0.080 ;
      RECT 1.000 -0.080 1.090 0.122 ;
      RECT 0.734 -0.080 1.000 0.080 ;
      RECT 0.644 -0.080 0.734 0.122 ;
      RECT 0.306 -0.080 0.644 0.080 ;
      RECT 0.216 -0.080 0.306 0.122 ;
      RECT 0.000 -0.080 0.216 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.250 1.120 1.400 1.280 ;
      RECT 1.160 0.971 1.250 1.280 ;
      RECT 0.335 1.120 1.160 1.280 ;
      RECT 0.245 1.065 0.335 1.280 ;
      RECT 0.000 1.120 0.245 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.181 0.301 1.242 0.760 ;
      RECT 0.773 0.424 1.181 0.479 ;
      RECT 1.144 0.679 1.181 0.760 ;
      RECT 0.860 0.542 0.951 0.624 ;
      RECT 0.797 0.569 0.860 0.624 ;
      RECT 0.736 0.569 0.797 0.744 ;
      RECT 0.683 0.424 0.773 0.514 ;
      RECT 0.263 0.689 0.736 0.744 ;
      RECT 0.202 0.292 0.263 0.744 ;
      RECT 0.138 0.292 0.202 0.346 ;
      RECT 0.138 0.669 0.202 0.744 ;
      RECT 0.048 0.265 0.138 0.346 ;
      RECT 0.048 0.669 0.138 0.750 ;
  END
END NOR4BBX1

MACRO NOR4BXL
  CLASS CORE ;
  FOREIGN NOR4BXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.036 0.439 1.040 0.494 ;
      RECT 0.972 0.287 1.036 0.801 ;
      RECT 0.889 0.287 0.972 0.342 ;
      RECT 0.917 0.720 0.972 0.801 ;
      RECT 0.428 0.261 0.889 0.342 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.336 0.556 0.400 0.755 ;
      RECT 0.307 0.700 0.336 0.755 ;
      RECT 0.243 0.700 0.307 0.761 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.528 0.557 0.603 0.638 ;
      RECT 0.508 0.439 0.528 0.638 ;
      RECT 0.464 0.439 0.508 0.612 ;
      RECT 0.426 0.439 0.464 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.697 0.413 0.878 0.513 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.395 0.144 0.532 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 -0.080 1.100 0.080 ;
      RECT 0.950 -0.080 1.044 0.122 ;
      RECT 0.678 -0.080 0.950 0.080 ;
      RECT 0.583 -0.080 0.678 0.122 ;
      RECT 0.328 -0.080 0.583 0.080 ;
      RECT 0.233 -0.080 0.328 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.300 1.120 1.100 1.280 ;
      RECT 0.206 1.078 0.300 1.280 ;
      RECT 0.000 1.120 0.206 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.731 0.594 0.908 0.649 ;
      RECT 0.667 0.594 0.731 0.876 ;
      RECT 0.144 0.821 0.667 0.876 ;
      RECT 0.208 0.273 0.272 0.643 ;
      RECT 0.144 0.273 0.208 0.327 ;
      RECT 0.144 0.588 0.208 0.643 ;
      RECT 0.050 0.244 0.144 0.327 ;
      RECT 0.081 0.588 0.144 0.876 ;
      RECT 0.050 0.720 0.081 0.801 ;
  END
END NOR4BXL

MACRO NOR4BX4
  CLASS CORE ;
  FOREIGN NOR4BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.142 0.567 3.162 0.900 ;
      RECT 3.080 0.282 3.142 0.923 ;
      RECT 2.908 0.282 3.080 0.337 ;
      RECT 3.060 0.567 3.080 0.923 ;
      RECT 2.393 0.868 3.060 0.923 ;
      RECT 2.816 0.256 2.908 0.337 ;
      RECT 2.516 0.282 2.816 0.337 ;
      RECT 2.424 0.256 2.516 0.337 ;
      RECT 0.916 0.282 2.424 0.337 ;
      RECT 2.364 0.867 2.393 0.948 ;
      RECT 2.302 0.867 2.364 1.008 ;
      RECT 1.030 0.954 2.302 1.008 ;
      RECT 0.939 0.954 1.030 1.035 ;
      RECT 0.824 0.256 0.916 0.337 ;
      RECT 0.528 0.282 0.824 0.337 ;
      RECT 0.436 0.256 0.528 0.337 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.970 0.429 3.007 0.510 ;
      RECT 2.908 0.429 2.970 0.758 ;
      RECT 1.720 0.704 2.908 0.758 ;
      RECT 1.705 0.704 1.720 0.761 ;
      RECT 1.675 0.618 1.705 0.761 ;
      RECT 1.613 0.618 1.675 0.899 ;
      RECT 0.409 0.844 1.613 0.899 ;
      RECT 0.347 0.526 0.409 0.899 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.789 0.476 2.819 0.573 ;
      RECT 2.727 0.476 2.789 0.648 ;
      RECT 1.945 0.593 2.727 0.648 ;
      RECT 1.883 0.502 1.945 0.648 ;
      RECT 1.853 0.502 1.883 0.583 ;
      RECT 1.815 0.502 1.853 0.573 ;
      RECT 1.479 0.502 1.815 0.557 ;
      RECT 1.449 0.502 1.479 0.583 ;
      RECT 1.385 0.502 1.449 0.789 ;
      RECT 1.302 0.706 1.385 0.789 ;
      RECT 0.605 0.735 1.302 0.789 ;
      RECT 0.528 0.556 0.605 0.789 ;
      RECT 0.513 0.556 0.528 0.637 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.547 0.457 2.638 0.538 ;
      RECT 2.191 0.483 2.547 0.538 ;
      RECT 2.117 0.433 2.191 0.538 ;
      RECT 2.055 0.392 2.117 0.538 ;
      RECT 1.277 0.392 2.055 0.446 ;
      RECT 1.215 0.392 1.277 0.637 ;
      RECT 1.185 0.556 1.215 0.637 ;
      RECT 0.785 0.573 1.185 0.627 ;
      RECT 0.694 0.563 0.785 0.644 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.046 0.439 0.137 0.608 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.106 -0.080 3.200 0.080 ;
      RECT 3.014 -0.080 3.106 0.212 ;
      RECT 2.711 -0.080 3.014 0.080 ;
      RECT 2.620 -0.080 2.711 0.212 ;
      RECT 2.322 -0.080 2.620 0.080 ;
      RECT 2.230 -0.080 2.322 0.212 ;
      RECT 1.114 -0.080 2.230 0.080 ;
      RECT 1.022 -0.080 1.114 0.212 ;
      RECT 0.722 -0.080 1.022 0.080 ;
      RECT 0.630 -0.080 0.722 0.211 ;
      RECT 0.334 -0.080 0.630 0.080 ;
      RECT 0.242 -0.080 0.334 0.211 ;
      RECT 0.000 -0.080 0.242 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.106 1.120 3.200 1.280 ;
      RECT 3.014 1.078 3.106 1.280 ;
      RECT 1.712 1.120 3.014 1.280 ;
      RECT 1.620 1.078 1.712 1.280 ;
      RECT 0.349 1.120 1.620 1.280 ;
      RECT 0.257 1.078 0.349 1.280 ;
      RECT 0.000 1.120 0.257 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.951 0.415 1.042 0.510 ;
      RECT 0.281 0.415 0.951 0.470 ;
      RECT 0.220 0.320 0.281 0.869 ;
      RECT 0.140 0.320 0.220 0.375 ;
      RECT 0.140 0.814 0.220 0.869 ;
      RECT 0.048 0.224 0.140 0.375 ;
      RECT 0.048 0.814 0.140 0.895 ;
  END
END NOR4BX4

MACRO NOR4BX2
  CLASS CORE ;
  FOREIGN NOR4BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.675 0.192 1.737 0.894 ;
      RECT 1.658 0.192 1.675 0.306 ;
      RECT 1.140 0.839 1.675 0.894 ;
      RECT 0.949 0.192 1.658 0.246 ;
      RECT 1.058 0.833 1.140 0.900 ;
      RECT 0.965 0.826 1.058 0.907 ;
      RECT 0.856 0.179 0.949 0.260 ;
      RECT 0.442 0.192 0.856 0.246 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.580 0.557 1.612 0.638 ;
      RECT 1.519 0.557 1.580 0.761 ;
      RECT 1.518 0.570 1.519 0.761 ;
      RECT 0.419 0.706 1.518 0.761 ;
      RECT 0.390 0.700 0.419 0.761 ;
      RECT 0.297 0.569 0.390 0.761 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.396 1.561 0.500 ;
      RECT 1.400 0.343 1.480 0.500 ;
      RECT 0.682 0.343 1.400 0.398 ;
      RECT 0.641 0.343 0.682 0.439 ;
      RECT 0.578 0.343 0.641 0.533 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.139 0.452 1.276 0.627 ;
      RECT 0.840 0.452 1.139 0.507 ;
      RECT 0.747 0.452 0.840 0.533 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.433 0.322 0.513 ;
      RECT 0.160 0.395 0.222 0.513 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.156 -0.080 1.800 0.080 ;
      RECT 1.064 -0.080 1.156 0.122 ;
      RECT 0.742 -0.080 1.064 0.080 ;
      RECT 0.649 -0.080 0.742 0.122 ;
      RECT 0.338 -0.080 0.649 0.080 ;
      RECT 0.245 -0.080 0.338 0.198 ;
      RECT 0.000 -0.080 0.245 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.724 1.120 1.800 1.280 ;
      RECT 1.631 1.078 1.724 1.280 ;
      RECT 0.327 1.120 1.631 1.280 ;
      RECT 0.235 1.078 0.327 1.280 ;
      RECT 0.000 1.120 0.235 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.926 0.570 1.023 0.643 ;
      RECT 0.515 0.588 0.926 0.643 ;
      RECT 0.453 0.301 0.515 0.643 ;
      RECT 0.359 0.301 0.453 0.356 ;
      RECT 0.296 0.268 0.359 0.356 ;
      RECT 0.142 0.268 0.296 0.323 ;
      RECT 0.097 0.217 0.142 0.323 ;
      RECT 0.097 0.683 0.142 0.876 ;
      RECT 0.034 0.217 0.097 0.876 ;
  END
END NOR4BX2

MACRO NOR4BX1
  CLASS CORE ;
  FOREIGN NOR4BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.036 0.439 1.040 0.494 ;
      RECT 0.972 0.288 1.036 0.799 ;
      RECT 0.889 0.288 0.972 0.343 ;
      RECT 0.917 0.718 0.972 0.799 ;
      RECT 0.428 0.262 0.889 0.343 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.336 0.556 0.400 0.755 ;
      RECT 0.307 0.700 0.336 0.755 ;
      RECT 0.243 0.700 0.307 0.761 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.528 0.557 0.603 0.638 ;
      RECT 0.508 0.439 0.528 0.638 ;
      RECT 0.464 0.439 0.508 0.612 ;
      RECT 0.426 0.439 0.464 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.697 0.413 0.878 0.513 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.143 0.395 0.144 0.531 ;
      RECT 0.049 0.395 0.143 0.532 ;
      RECT 0.038 0.395 0.049 0.531 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 -0.080 1.100 0.080 ;
      RECT 0.950 -0.080 1.044 0.122 ;
      RECT 0.678 -0.080 0.950 0.080 ;
      RECT 0.583 -0.080 0.678 0.122 ;
      RECT 0.328 -0.080 0.583 0.080 ;
      RECT 0.233 -0.080 0.328 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.328 1.120 1.100 1.280 ;
      RECT 0.233 1.078 0.328 1.280 ;
      RECT 0.000 1.120 0.233 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.731 0.594 0.908 0.649 ;
      RECT 0.667 0.594 0.731 0.876 ;
      RECT 0.144 0.821 0.667 0.876 ;
      RECT 0.208 0.273 0.272 0.643 ;
      RECT 0.144 0.273 0.208 0.327 ;
      RECT 0.144 0.588 0.208 0.643 ;
      RECT 0.050 0.246 0.144 0.327 ;
      RECT 0.081 0.588 0.144 0.876 ;
      RECT 0.050 0.707 0.081 0.788 ;
  END
END NOR4BX1

MACRO NOR4X2
  CLASS CORE ;
  FOREIGN NOR4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.287 1.542 1.008 ;
      RECT 0.813 0.287 1.480 0.342 ;
      RECT 1.460 0.894 1.480 1.008 ;
      RECT 0.853 0.954 1.460 1.008 ;
      RECT 0.761 0.954 0.853 1.035 ;
      RECT 0.722 0.261 0.813 0.342 ;
      RECT 0.338 0.287 0.722 0.342 ;
      RECT 0.246 0.261 0.338 0.342 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.387 0.556 1.417 0.637 ;
      RECT 1.325 0.556 1.387 0.899 ;
      RECT 0.238 0.844 1.325 0.899 ;
      RECT 0.176 0.556 0.238 0.899 ;
      RECT 0.055 0.556 0.176 0.637 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.174 0.396 1.236 0.789 ;
      RECT 1.145 0.396 1.174 0.477 ;
      RECT 0.475 0.735 1.174 0.789 ;
      RECT 0.427 0.706 0.475 0.789 ;
      RECT 0.365 0.556 0.427 0.789 ;
      RECT 0.335 0.556 0.365 0.637 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.069 0.556 1.099 0.637 ;
      RECT 1.007 0.444 1.069 0.637 ;
      RECT 0.653 0.444 1.007 0.499 ;
      RECT 0.607 0.439 0.653 0.499 ;
      RECT 0.517 0.439 0.607 0.538 ;
      RECT 0.516 0.457 0.517 0.538 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.710 0.555 0.878 0.636 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.018 -0.080 1.600 0.080 ;
      RECT 0.927 -0.080 1.018 0.122 ;
      RECT 0.593 -0.080 0.927 0.080 ;
      RECT 0.501 -0.080 0.593 0.122 ;
      RECT 0.140 -0.080 0.501 0.080 ;
      RECT 0.048 -0.080 0.140 0.225 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.534 1.120 1.600 1.280 ;
      RECT 1.442 1.078 1.534 1.280 ;
      RECT 0.140 1.120 1.442 1.280 ;
      RECT 0.048 1.078 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
END NOR4X2

MACRO NOR4X1
  CLASS CORE ;
  FOREIGN NOR4X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.976 0.269 1.040 0.761 ;
      RECT 0.261 0.269 0.976 0.350 ;
      RECT 0.879 0.706 0.976 0.761 ;
      RECT 0.785 0.698 0.879 0.890 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.156 0.542 0.157 0.623 ;
      RECT 0.062 0.542 0.156 0.700 ;
      RECT 0.057 0.573 0.062 0.627 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.243 0.421 0.440 0.519 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.593 0.433 0.626 0.514 ;
      RECT 0.529 0.433 0.593 0.761 ;
      RECT 0.426 0.700 0.529 0.761 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.811 0.420 0.906 0.560 ;
      RECT 0.793 0.439 0.811 0.494 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 -0.080 1.100 0.080 ;
      RECT 0.956 -0.080 1.050 0.122 ;
      RECT 0.611 -0.080 0.956 0.080 ;
      RECT 0.517 -0.080 0.611 0.122 ;
      RECT 0.144 -0.080 0.517 0.080 ;
      RECT 0.050 -0.080 0.144 0.122 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.144 1.120 1.100 1.280 ;
      RECT 0.050 1.078 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
END NOR4X1

MACRO NOR3BX4
  CLASS CORE ;
  FOREIGN NOR3BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.920 0.433 1.961 0.852 ;
      RECT 1.857 0.268 1.920 0.852 ;
      RECT 1.431 0.268 1.857 0.323 ;
      RECT 1.807 0.771 1.857 0.852 ;
      RECT 1.052 0.771 1.807 0.826 ;
      RECT 1.368 0.165 1.431 0.323 ;
      RECT 1.337 0.165 1.368 0.246 ;
      RECT 1.011 0.192 1.337 0.246 ;
      RECT 1.032 0.771 1.052 0.839 ;
      RECT 0.968 0.771 1.032 0.867 ;
      RECT 0.917 0.165 1.011 0.246 ;
      RECT 0.876 0.812 0.968 0.867 ;
      RECT 0.592 0.192 0.917 0.246 ;
      RECT 0.782 0.812 0.876 0.893 ;
      RECT 0.499 0.165 0.592 0.246 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.295 0.414 1.455 0.495 ;
      RECT 1.231 0.301 1.295 0.495 ;
      RECT 0.486 0.301 1.231 0.356 ;
      RECT 0.423 0.301 0.486 0.627 ;
      RECT 0.366 0.536 0.423 0.617 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.561 0.523 1.624 0.606 ;
      RECT 1.128 0.551 1.561 0.606 ;
      RECT 1.098 0.520 1.128 0.606 ;
      RECT 1.034 0.411 1.098 0.606 ;
      RECT 1.032 0.411 1.034 0.500 ;
      RECT 0.668 0.411 1.032 0.465 ;
      RECT 0.658 0.411 0.668 0.513 ;
      RECT 0.565 0.411 0.658 0.514 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.284 0.306 0.304 0.361 ;
      RECT 0.220 0.306 0.284 0.519 ;
      RECT 0.180 0.438 0.220 0.519 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.629 -0.080 2.000 0.080 ;
      RECT 1.536 -0.080 1.629 0.198 ;
      RECT 1.222 -0.080 1.536 0.080 ;
      RECT 1.128 -0.080 1.222 0.122 ;
      RECT 0.802 -0.080 1.128 0.080 ;
      RECT 0.708 -0.080 0.802 0.122 ;
      RECT 0.394 -0.080 0.708 0.080 ;
      RECT 0.300 -0.080 0.394 0.198 ;
      RECT 0.000 -0.080 0.300 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.388 1.120 2.000 1.280 ;
      RECT 1.295 0.911 1.388 1.280 ;
      RECT 0.358 1.120 1.295 1.280 ;
      RECT 0.264 0.866 0.358 1.280 ;
      RECT 0.000 1.120 0.264 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.687 0.377 1.769 0.715 ;
      RECT 1.667 0.377 1.687 0.437 ;
      RECT 0.879 0.661 1.687 0.715 ;
      RECT 0.780 0.520 0.879 0.756 ;
      RECT 0.143 0.701 0.780 0.756 ;
      RECT 0.113 0.198 0.157 0.282 ;
      RECT 0.113 0.701 0.143 0.790 ;
      RECT 0.050 0.198 0.113 0.790 ;
  END
END NOR3BX4

MACRO NOR3BX2
  CLASS CORE ;
  FOREIGN NOR3BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.270 0.192 1.331 0.861 ;
      RECT 1.262 0.192 1.270 0.306 ;
      RECT 1.262 0.761 1.270 0.861 ;
      RECT 0.973 0.192 1.262 0.246 ;
      RECT 0.993 0.806 1.262 0.861 ;
      RECT 0.932 0.806 0.993 0.894 ;
      RECT 0.883 0.165 0.973 0.246 ;
      RECT 0.843 0.806 0.932 0.861 ;
      RECT 0.570 0.192 0.883 0.246 ;
      RECT 0.753 0.806 0.843 0.895 ;
      RECT 0.480 0.165 0.570 0.246 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.180 0.394 1.209 0.475 ;
      RECT 1.119 0.324 1.180 0.475 ;
      RECT 0.467 0.324 1.119 0.379 ;
      RECT 0.467 0.573 0.468 0.627 ;
      RECT 0.406 0.324 0.467 0.627 ;
      RECT 0.387 0.494 0.406 0.627 ;
      RECT 0.365 0.536 0.387 0.627 ;
      RECT 0.335 0.536 0.365 0.617 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.057 0.555 1.086 0.636 ;
      RECT 0.996 0.461 1.057 0.636 ;
      RECT 0.643 0.461 0.996 0.515 ;
      RECT 0.619 0.439 0.643 0.515 ;
      RECT 0.558 0.439 0.619 0.542 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.273 0.306 0.293 0.361 ;
      RECT 0.212 0.306 0.273 0.457 ;
      RECT 0.174 0.376 0.212 0.457 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.772 -0.080 1.400 0.080 ;
      RECT 0.681 -0.080 0.772 0.122 ;
      RECT 0.379 -0.080 0.681 0.080 ;
      RECT 0.289 -0.080 0.379 0.198 ;
      RECT 0.000 -0.080 0.289 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 1.120 1.400 1.280 ;
      RECT 1.246 0.932 1.336 1.280 ;
      RECT 0.345 1.120 1.246 1.280 ;
      RECT 0.255 0.897 0.345 1.280 ;
      RECT 0.000 1.120 0.255 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.846 0.570 0.875 0.625 ;
      RECT 0.785 0.570 0.846 0.751 ;
      RECT 0.138 0.696 0.785 0.751 ;
      RECT 0.109 0.198 0.151 0.282 ;
      RECT 0.109 0.670 0.138 0.751 ;
      RECT 0.048 0.198 0.109 0.751 ;
  END
END NOR3BX2

MACRO NOR3BX1
  CLASS CORE ;
  FOREIGN NOR3BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.003 0.269 1.067 0.894 ;
      RECT 0.486 0.269 1.003 0.350 ;
      RECT 0.878 0.839 1.003 0.894 ;
      RECT 0.783 0.839 0.878 0.924 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.489 0.573 0.490 0.627 ;
      RECT 0.307 0.536 0.489 0.627 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.553 0.414 0.756 0.511 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.286 0.306 0.307 0.361 ;
      RECT 0.222 0.306 0.286 0.457 ;
      RECT 0.182 0.376 0.222 0.457 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.792 -0.080 1.100 0.080 ;
      RECT 0.697 -0.080 0.792 0.122 ;
      RECT 0.415 -0.080 0.697 0.080 ;
      RECT 0.321 -0.080 0.415 0.122 ;
      RECT 0.000 -0.080 0.321 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.361 1.120 1.100 1.280 ;
      RECT 0.267 0.897 0.361 1.280 ;
      RECT 0.000 1.120 0.267 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.886 0.536 0.917 0.617 ;
      RECT 0.822 0.536 0.886 0.751 ;
      RECT 0.144 0.696 0.822 0.751 ;
      RECT 0.114 0.237 0.150 0.321 ;
      RECT 0.114 0.670 0.144 0.751 ;
      RECT 0.050 0.237 0.114 0.751 ;
  END
END NOR3BX1

MACRO NOR3X4
  CLASS CORE ;
  FOREIGN NOR3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.721 0.567 1.762 0.900 ;
      RECT 1.658 0.268 1.721 0.900 ;
      RECT 1.124 0.268 1.658 0.323 ;
      RECT 1.561 0.810 1.658 0.892 ;
      RECT 0.665 0.837 1.561 0.892 ;
      RECT 1.031 0.242 1.124 0.323 ;
      RECT 0.731 0.268 1.031 0.323 ;
      RECT 0.638 0.242 0.731 0.323 ;
      RECT 0.573 0.837 0.665 0.918 ;
      RECT 0.338 0.268 0.638 0.323 ;
      RECT 0.245 0.242 0.338 0.323 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.092 0.598 1.189 0.774 ;
      RECT 1.021 0.700 1.092 0.774 ;
      RECT 0.153 0.719 1.021 0.774 ;
      RECT 0.090 0.526 0.153 0.774 ;
      RECT 0.056 0.526 0.090 0.627 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.971 0.488 1.390 0.543 ;
      RECT 0.908 0.488 0.971 0.610 ;
      RECT 0.404 0.555 0.908 0.610 ;
      RECT 0.374 0.507 0.404 0.610 ;
      RECT 0.311 0.439 0.374 0.610 ;
      RECT 0.239 0.439 0.311 0.494 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.553 0.581 1.582 0.662 ;
      RECT 1.490 0.379 1.553 0.662 ;
      RECT 0.731 0.379 1.490 0.433 ;
      RECT 1.489 0.581 1.490 0.662 ;
      RECT 0.638 0.379 0.731 0.496 ;
      RECT 0.599 0.429 0.638 0.494 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.320 -0.080 1.800 0.080 ;
      RECT 1.227 -0.080 1.320 0.198 ;
      RECT 0.927 -0.080 1.227 0.080 ;
      RECT 0.835 -0.080 0.927 0.198 ;
      RECT 0.535 -0.080 0.835 0.080 ;
      RECT 0.442 -0.080 0.535 0.198 ;
      RECT 0.142 -0.080 0.442 0.080 ;
      RECT 0.049 -0.080 0.142 0.211 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.181 1.120 1.800 1.280 ;
      RECT 1.088 0.989 1.181 1.280 ;
      RECT 0.142 1.120 1.088 1.280 ;
      RECT 0.049 0.929 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
END NOR3X4

MACRO NOR3X2
  CLASS CORE ;
  FOREIGN NOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.255 1.240 0.855 ;
      RECT 0.754 0.255 1.175 0.310 ;
      RECT 1.154 0.767 1.175 0.855 ;
      RECT 0.687 0.800 1.154 0.855 ;
      RECT 0.658 0.151 0.754 0.344 ;
      RECT 0.591 0.800 0.687 0.890 ;
      RECT 0.349 0.289 0.658 0.344 ;
      RECT 0.253 0.151 0.349 0.344 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.007 0.537 1.088 0.744 ;
      RECT 0.214 0.689 1.007 0.744 ;
      RECT 0.149 0.573 0.214 0.744 ;
      RECT 0.118 0.573 0.149 0.707 ;
      RECT 0.058 0.573 0.118 0.627 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.913 0.377 0.943 0.458 ;
      RECT 0.848 0.377 0.913 0.635 ;
      RECT 0.847 0.377 0.848 0.458 ;
      RECT 0.416 0.580 0.848 0.635 ;
      RECT 0.415 0.458 0.416 0.635 ;
      RECT 0.352 0.445 0.415 0.635 ;
      RECT 0.321 0.445 0.352 0.539 ;
      RECT 0.311 0.445 0.321 0.500 ;
      RECT 0.246 0.439 0.311 0.500 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.498 0.439 0.682 0.525 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.552 -0.080 1.300 0.080 ;
      RECT 0.456 -0.080 0.552 0.211 ;
      RECT 0.146 -0.080 0.456 0.080 ;
      RECT 0.051 -0.080 0.146 0.211 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 1.120 1.300 1.280 ;
      RECT 1.109 0.925 1.204 1.280 ;
      RECT 0.146 1.120 1.109 1.280 ;
      RECT 0.051 0.876 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
END NOR3X2

MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.666 0.269 0.668 0.894 ;
      RECT 0.607 0.269 0.666 0.924 ;
      RECT 0.196 0.269 0.607 0.350 ;
      RECT 0.557 0.839 0.607 0.924 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.137 0.536 0.138 0.617 ;
      RECT 0.048 0.536 0.137 0.694 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.421 0.361 0.561 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.517 0.536 0.546 0.617 ;
      RECT 0.456 0.536 0.517 0.761 ;
      RECT 0.407 0.706 0.456 0.761 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 -0.080 0.700 0.080 ;
      RECT 0.345 -0.080 0.435 0.122 ;
      RECT 0.138 -0.080 0.345 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.138 1.120 0.700 1.280 ;
      RECT 0.048 0.900 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
END NOR3X1

MACRO NOR2BXL
  CLASS CORE ;
  FOREIGN NOR2BXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.605 0.295 0.666 0.798 ;
      RECT 0.501 0.295 0.605 0.350 ;
      RECT 0.562 0.706 0.605 0.798 ;
      RECT 0.411 0.269 0.501 0.350 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.411 0.567 0.525 0.633 ;
      RECT 0.321 0.567 0.411 0.662 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.433 0.138 0.581 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 -0.080 0.700 0.080 ;
      RECT 0.562 -0.080 0.652 0.122 ;
      RECT 0.313 -0.080 0.562 0.080 ;
      RECT 0.223 -0.080 0.313 0.122 ;
      RECT 0.000 -0.080 0.223 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.302 1.120 0.700 1.280 ;
      RECT 0.212 1.078 0.302 1.280 ;
      RECT 0.000 1.120 0.212 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.260 0.421 0.544 0.502 ;
      RECT 0.199 0.321 0.260 0.762 ;
      RECT 0.138 0.321 0.199 0.376 ;
      RECT 0.138 0.707 0.199 0.762 ;
      RECT 0.048 0.295 0.138 0.376 ;
      RECT 0.048 0.707 0.138 0.788 ;
  END
END NOR2BXL

MACRO NOR2BX4
  CLASS CORE ;
  FOREIGN NOR2BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.262 0.264 1.363 0.786 ;
      RECT 0.973 0.264 1.262 0.336 ;
      RECT 1.252 0.693 1.262 0.786 ;
      RECT 0.573 0.705 1.252 0.786 ;
      RECT 0.883 0.255 0.973 0.336 ;
      RECT 0.570 0.281 0.883 0.336 ;
      RECT 0.480 0.255 0.570 0.336 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.936 0.563 1.026 0.650 ;
      RECT 0.468 0.595 0.936 0.650 ;
      RECT 0.411 0.565 0.468 0.650 ;
      RECT 0.321 0.521 0.411 0.650 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.034 0.436 0.138 0.571 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.177 -0.080 1.400 0.080 ;
      RECT 1.087 -0.080 1.177 0.122 ;
      RECT 0.772 -0.080 1.087 0.080 ;
      RECT 0.681 -0.080 0.772 0.122 ;
      RECT 0.366 -0.080 0.681 0.080 ;
      RECT 0.276 -0.080 0.366 0.122 ;
      RECT 0.000 -0.080 0.276 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.013 1.120 1.400 1.280 ;
      RECT 0.923 1.078 1.013 1.280 ;
      RECT 0.313 1.117 0.923 1.280 ;
      RECT 0.223 1.078 0.313 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.139 0.392 1.200 0.546 ;
      RECT 0.668 0.392 1.139 0.446 ;
      RECT 0.578 0.392 0.668 0.538 ;
      RECT 0.260 0.392 0.578 0.446 ;
      RECT 0.199 0.307 0.260 0.848 ;
      RECT 0.164 0.307 0.199 0.362 ;
      RECT 0.138 0.793 0.199 0.848 ;
      RECT 0.074 0.281 0.164 0.362 ;
      RECT 0.048 0.793 0.138 0.874 ;
  END
END NOR2BX4

MACRO NOR2BX2
  CLASS CORE ;
  FOREIGN NOR2BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.997 0.308 1.061 0.767 ;
      RECT 0.850 0.308 0.997 0.363 ;
      RECT 0.976 0.706 0.997 0.767 ;
      RECT 0.689 0.712 0.976 0.767 ;
      RECT 0.756 0.282 0.850 0.363 ;
      RECT 0.594 0.712 0.689 0.793 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.847 0.418 0.928 0.565 ;
      RECT 0.511 0.418 0.847 0.473 ;
      RECT 0.436 0.300 0.511 0.473 ;
      RECT 0.406 0.300 0.436 0.514 ;
      RECT 0.357 0.418 0.406 0.514 ;
      RECT 0.342 0.433 0.357 0.514 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.050 0.457 0.144 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 -0.080 1.100 0.080 ;
      RECT 0.956 -0.080 1.050 0.228 ;
      RECT 0.636 -0.080 0.956 0.080 ;
      RECT 0.542 -0.080 0.636 0.122 ;
      RECT 0.000 -0.080 0.542 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 1.120 1.100 1.280 ;
      RECT 0.956 1.078 1.050 1.280 ;
      RECT 0.322 1.120 0.956 1.280 ;
      RECT 0.228 1.078 0.322 1.280 ;
      RECT 0.000 1.120 0.228 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.622 0.538 0.717 0.626 ;
      RECT 0.272 0.571 0.622 0.626 ;
      RECT 0.208 0.312 0.272 0.802 ;
      RECT 0.144 0.312 0.208 0.367 ;
      RECT 0.144 0.748 0.208 0.802 ;
      RECT 0.050 0.286 0.144 0.367 ;
      RECT 0.050 0.748 0.144 0.829 ;
  END
END NOR2BX2

MACRO NOR2BX1
  CLASS CORE ;
  FOREIGN NOR2BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.605 0.295 0.666 0.858 ;
      RECT 0.501 0.295 0.605 0.350 ;
      RECT 0.562 0.706 0.605 0.858 ;
      RECT 0.411 0.269 0.501 0.350 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.411 0.567 0.525 0.633 ;
      RECT 0.321 0.567 0.411 0.670 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.486 0.138 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 -0.080 0.700 0.080 ;
      RECT 0.562 -0.080 0.652 0.122 ;
      RECT 0.353 -0.080 0.562 0.080 ;
      RECT 0.263 -0.080 0.353 0.122 ;
      RECT 0.000 -0.080 0.263 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.302 1.120 0.700 1.280 ;
      RECT 0.212 0.916 0.302 1.280 ;
      RECT 0.000 1.120 0.212 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.461 0.430 0.544 0.511 ;
      RECT 0.260 0.443 0.461 0.498 ;
      RECT 0.199 0.323 0.260 0.770 ;
      RECT 0.138 0.323 0.199 0.385 ;
      RECT 0.138 0.715 0.199 0.770 ;
      RECT 0.048 0.304 0.138 0.385 ;
      RECT 0.048 0.715 0.138 0.796 ;
  END
END NOR2BX1

MACRO NOR2XL
  CLASS CORE ;
  FOREIGN NOR2XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.491 0.295 0.561 0.774 ;
      RECT 0.352 0.295 0.491 0.350 ;
      RECT 0.442 0.626 0.491 0.774 ;
      RECT 0.248 0.269 0.352 0.350 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.164 0.567 0.255 0.633 ;
      RECT 0.061 0.548 0.164 0.633 ;
      RECT 0.042 0.567 0.061 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.242 0.406 0.421 0.502 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.545 -0.080 0.600 0.080 ;
      RECT 0.442 -0.080 0.545 0.122 ;
      RECT 0.158 -0.080 0.442 0.080 ;
      RECT 0.055 -0.080 0.158 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 1.120 0.600 1.280 ;
      RECT 0.055 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.055 1.280 ;
     END
  END VDD
END NOR2XL

MACRO NOR2X4
  CLASS CORE ;
  FOREIGN NOR2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 0.433 1.261 0.767 ;
      RECT 1.244 0.265 1.249 0.767 ;
      RECT 1.165 0.265 1.244 0.840 ;
      RECT 0.765 0.265 1.165 0.337 ;
      RECT 1.154 0.433 1.165 0.840 ;
      RECT 1.148 0.693 1.154 0.840 ;
      RECT 0.428 0.760 1.148 0.840 ;
      RECT 0.670 0.256 0.765 0.337 ;
      RECT 0.360 0.282 0.670 0.337 ;
      RECT 0.265 0.256 0.360 0.337 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.827 0.561 0.858 0.642 ;
      RECT 0.763 0.561 0.827 0.705 ;
      RECT 0.311 0.650 0.763 0.705 ;
      RECT 0.246 0.650 0.311 0.761 ;
      RECT 0.234 0.650 0.246 0.707 ;
      RECT 0.169 0.492 0.234 0.707 ;
      RECT 0.138 0.492 0.169 0.573 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.055 0.464 1.086 0.545 ;
      RECT 0.990 0.394 1.055 0.545 ;
      RECT 0.523 0.394 0.990 0.449 ;
      RECT 0.459 0.394 0.523 0.525 ;
      RECT 0.432 0.439 0.459 0.525 ;
      RECT 0.428 0.470 0.432 0.525 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.979 -0.080 1.300 0.080 ;
      RECT 0.884 -0.080 0.979 0.122 ;
      RECT 0.563 -0.080 0.884 0.080 ;
      RECT 0.467 -0.080 0.563 0.211 ;
      RECT 0.146 -0.080 0.467 0.080 ;
      RECT 0.051 -0.080 0.146 0.298 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.895 1.120 1.300 1.280 ;
      RECT 0.799 1.078 0.895 1.280 ;
      RECT 0.152 1.120 0.799 1.280 ;
      RECT 0.056 1.078 0.152 1.280 ;
      RECT 0.000 1.120 0.056 1.280 ;
     END
  END VDD
END NOR2X4

MACRO NOR2X2
  CLASS CORE ;
  FOREIGN NOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.862 0.308 0.867 0.761 ;
      RECT 0.805 0.308 0.862 0.767 ;
      RECT 0.655 0.308 0.805 0.363 ;
      RECT 0.779 0.706 0.805 0.767 ;
      RECT 0.496 0.712 0.779 0.767 ;
      RECT 0.562 0.170 0.655 0.363 ;
      RECT 0.404 0.712 0.496 0.793 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 0.418 0.742 0.564 ;
      RECT 0.229 0.418 0.652 0.473 ;
      RECT 0.120 0.418 0.229 0.518 ;
      RECT 0.059 0.418 0.120 0.494 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.327 0.538 0.502 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.228 ;
      RECT 0.458 -0.080 0.758 0.080 ;
      RECT 0.365 -0.080 0.458 0.340 ;
      RECT 0.000 -0.080 0.365 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.758 1.078 0.851 1.280 ;
      RECT 0.142 1.120 0.758 1.280 ;
      RECT 0.049 1.078 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
END NOR2X2

MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.491 0.295 0.561 0.774 ;
      RECT 0.352 0.295 0.491 0.350 ;
      RECT 0.442 0.626 0.491 0.774 ;
      RECT 0.248 0.269 0.352 0.350 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.164 0.567 0.255 0.643 ;
      RECT 0.061 0.548 0.164 0.643 ;
      RECT 0.042 0.567 0.061 0.643 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.242 0.407 0.421 0.502 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.545 -0.080 0.600 0.080 ;
      RECT 0.442 -0.080 0.545 0.122 ;
      RECT 0.158 -0.080 0.442 0.080 ;
      RECT 0.055 -0.080 0.158 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 1.120 0.600 1.280 ;
      RECT 0.055 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.055 1.280 ;
     END
  END VDD
END NOR2X1

MACRO NAND4BBX1
  CLASS CORE ;
  FOREIGN NAND4BBX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.343 0.573 1.367 0.933 ;
      RECT 1.306 0.201 1.343 0.933 ;
      RECT 1.282 0.201 1.306 0.627 ;
      RECT 0.878 0.879 1.306 0.933 ;
      RECT 1.262 0.201 1.282 0.306 ;
      RECT 0.964 0.201 1.262 0.256 ;
      RECT 0.874 0.201 0.964 0.282 ;
      RECT 0.817 0.742 0.878 0.933 ;
      RECT 0.788 0.742 0.817 0.839 ;
      RECT 0.737 0.755 0.788 0.839 ;
      RECT 0.582 0.755 0.737 0.810 ;
      RECT 0.517 0.742 0.582 0.810 ;
      RECT 0.427 0.742 0.517 0.823 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.412 0.439 0.468 0.494 ;
      RECT 0.351 0.439 0.412 0.600 ;
      RECT 0.327 0.519 0.351 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.610 0.439 0.643 0.494 ;
      RECT 0.549 0.439 0.610 0.636 ;
      RECT 0.502 0.555 0.549 0.636 ;
     END
  END C

  PIN BN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.041 0.433 0.142 0.574 ;
     END
  END BN

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.188 0.498 1.201 0.579 ;
      RECT 1.070 0.498 1.188 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.352 -0.080 1.400 0.080 ;
      RECT 1.262 -0.080 1.352 0.122 ;
      RECT 0.316 -0.080 1.262 0.080 ;
      RECT 0.098 -0.080 0.316 0.122 ;
      RECT 0.000 -0.080 0.098 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.077 1.120 1.400 1.280 ;
      RECT 0.957 1.078 1.077 1.280 ;
      RECT 0.697 1.120 0.957 1.280 ;
      RECT 0.607 1.078 0.697 1.280 ;
      RECT 0.337 1.120 0.607 1.280 ;
      RECT 0.322 1.078 0.337 1.280 ;
      RECT 0.261 1.065 0.322 1.280 ;
      RECT 0.247 1.078 0.261 1.280 ;
      RECT 0.000 1.120 0.247 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.005 0.755 1.245 0.810 ;
      RECT 1.059 0.311 1.149 0.392 ;
      RECT 1.005 0.337 1.059 0.392 ;
      RECT 0.944 0.337 1.005 0.810 ;
      RECT 0.890 0.419 0.944 0.500 ;
      RECT 0.738 0.302 0.799 0.636 ;
      RECT 0.264 0.302 0.738 0.357 ;
      RECT 0.709 0.555 0.738 0.636 ;
      RECT 0.203 0.302 0.264 0.801 ;
      RECT 0.138 0.302 0.203 0.357 ;
      RECT 0.138 0.746 0.203 0.801 ;
      RECT 0.048 0.293 0.138 0.374 ;
      RECT 0.048 0.746 0.138 0.827 ;
  END
END NAND4BBX1

MACRO NAND4BXL
  CLASS CORE ;
  FOREIGN NAND4BXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.668 0.839 0.857 0.894 ;
      RECT 0.672 0.252 0.767 0.333 ;
      RECT 0.639 0.279 0.672 0.333 ;
      RECT 0.639 0.839 0.668 0.939 ;
      RECT 0.575 0.279 0.639 0.939 ;
      RECT 0.490 0.858 0.575 0.939 ;
      RECT 0.300 0.885 0.490 0.939 ;
      RECT 0.206 0.858 0.300 0.939 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.078 0.439 0.167 0.600 ;
      RECT 0.060 0.439 0.078 0.599 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.661 0.383 0.767 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.368 0.433 0.511 0.532 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.874 0.546 1.061 0.652 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.957 -0.080 1.100 0.080 ;
      RECT 0.863 -0.080 0.957 0.122 ;
      RECT 0.144 -0.080 0.863 0.080 ;
      RECT 0.050 -0.080 0.144 0.122 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.882 1.120 1.100 1.280 ;
      RECT 0.787 1.078 0.882 1.280 ;
      RECT 0.511 1.120 0.787 1.280 ;
      RECT 0.417 1.078 0.511 1.280 ;
      RECT 0.144 1.120 0.417 1.280 ;
      RECT 0.050 1.078 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.007 0.806 1.037 0.887 ;
      RECT 0.943 0.724 1.007 0.887 ;
      RECT 0.960 0.320 0.990 0.401 ;
      RECT 0.896 0.320 0.960 0.482 ;
      RECT 0.769 0.724 0.943 0.779 ;
      RECT 0.769 0.427 0.896 0.482 ;
      RECT 0.706 0.427 0.769 0.779 ;
  END
END NAND4BXL

MACRO NAND4BX4
  CLASS CORE ;
  FOREIGN NAND4BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.983 0.567 2.985 0.900 ;
      RECT 2.974 0.288 2.983 0.900 ;
      RECT 2.921 0.288 2.974 0.942 ;
      RECT 2.316 0.288 2.921 0.343 ;
      RECT 2.882 0.567 2.921 0.942 ;
      RECT 2.294 0.870 2.882 0.942 ;
      RECT 2.225 0.150 2.316 0.343 ;
      RECT 0.467 0.870 2.294 0.937 ;
      RECT 1.002 0.207 2.225 0.274 ;
      RECT 0.910 0.150 1.002 0.343 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.815 0.426 2.859 0.507 ;
      RECT 2.769 0.426 2.815 0.815 ;
      RECT 2.753 0.439 2.769 0.815 ;
      RECT 1.659 0.761 2.753 0.815 ;
      RECT 1.568 0.735 1.659 0.815 ;
      RECT 0.475 0.761 1.568 0.815 ;
      RECT 0.453 0.706 0.475 0.815 ;
      RECT 0.413 0.519 0.453 0.815 ;
      RECT 0.391 0.519 0.413 0.761 ;
      RECT 0.361 0.519 0.391 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.668 0.519 2.683 0.600 ;
      RECT 2.591 0.519 2.668 0.633 ;
      RECT 2.589 0.573 2.591 0.633 ;
      RECT 2.547 0.573 2.589 0.706 ;
      RECT 2.527 0.579 2.547 0.706 ;
      RECT 1.916 0.651 2.527 0.706 ;
      RECT 1.825 0.625 1.916 0.706 ;
      RECT 1.401 0.625 1.825 0.680 ;
      RECT 1.309 0.625 1.401 0.706 ;
      RECT 0.653 0.651 1.309 0.706 ;
      RECT 0.591 0.519 0.653 0.706 ;
      RECT 0.544 0.519 0.591 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.451 0.515 2.465 0.596 ;
      RECT 2.349 0.433 2.451 0.596 ;
      RECT 2.104 0.542 2.349 0.596 ;
      RECT 2.003 0.510 2.104 0.596 ;
      RECT 1.222 0.510 2.003 0.564 ;
      RECT 1.121 0.510 1.222 0.596 ;
      RECT 0.824 0.542 1.121 0.596 ;
      RECT 0.723 0.515 0.824 0.596 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.144 0.574 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.974 -0.080 3.200 0.080 ;
      RECT 2.882 -0.080 2.974 0.122 ;
      RECT 1.659 -0.080 2.882 0.080 ;
      RECT 1.568 -0.080 1.659 0.122 ;
      RECT 0.345 -0.080 1.568 0.080 ;
      RECT 0.253 -0.080 0.345 0.122 ;
      RECT 0.000 -0.080 0.253 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.951 1.120 3.200 1.280 ;
      RECT 2.859 1.078 2.951 1.280 ;
      RECT 2.568 1.120 2.859 1.280 ;
      RECT 2.477 1.078 2.568 1.280 ;
      RECT 2.199 1.120 2.477 1.280 ;
      RECT 2.078 1.078 2.199 1.280 ;
      RECT 1.149 1.120 2.078 1.280 ;
      RECT 1.028 1.078 1.149 1.280 ;
      RECT 0.750 1.120 1.028 1.280 ;
      RECT 0.659 1.078 0.750 1.280 ;
      RECT 0.368 1.120 0.659 1.280 ;
      RECT 0.276 1.078 0.368 1.280 ;
      RECT 0.000 1.120 0.276 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.180 0.400 2.281 0.487 ;
      RECT 1.010 0.400 2.180 0.455 ;
      RECT 0.909 0.400 1.010 0.487 ;
      RECT 0.272 0.400 0.909 0.455 ;
      RECT 0.210 0.302 0.272 0.856 ;
      RECT 0.140 0.302 0.210 0.357 ;
      RECT 0.140 0.801 0.210 0.856 ;
      RECT 0.048 0.276 0.140 0.357 ;
      RECT 0.048 0.801 0.140 0.882 ;
  END
END NAND4BX4

MACRO NAND4BX2
  CLASS CORE ;
  FOREIGN NAND4BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.740 0.195 1.741 0.633 ;
      RECT 1.665 0.195 1.740 0.973 ;
      RECT 1.658 0.195 1.665 0.306 ;
      RECT 1.658 0.564 1.665 0.973 ;
      RECT 0.987 0.195 1.658 0.262 ;
      RECT 1.045 0.901 1.658 0.973 ;
      RECT 0.963 0.870 1.045 0.973 ;
      RECT 0.895 0.150 0.987 0.343 ;
      RECT 0.439 0.870 0.963 0.942 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.357 0.761 1.450 0.842 ;
      RECT 0.481 0.761 1.357 0.815 ;
      RECT 0.424 0.706 0.481 0.815 ;
      RECT 0.419 0.519 0.424 0.815 ;
      RECT 0.361 0.519 0.419 0.761 ;
      RECT 0.340 0.519 0.361 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.377 0.573 1.381 0.627 ;
      RECT 1.347 0.519 1.377 0.627 ;
      RECT 1.285 0.519 1.347 0.706 ;
      RECT 0.627 0.651 1.285 0.706 ;
      RECT 0.565 0.519 0.627 0.706 ;
      RECT 0.521 0.519 0.565 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.188 0.439 1.201 0.494 ;
      RECT 1.118 0.433 1.188 0.596 ;
      RECT 1.085 0.514 1.118 0.596 ;
      RECT 0.800 0.542 1.085 0.596 ;
      RECT 0.698 0.515 0.800 0.596 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.146 0.574 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.653 -0.080 1.800 0.080 ;
      RECT 1.560 -0.080 1.653 0.122 ;
      RECT 0.322 -0.080 1.560 0.080 ;
      RECT 0.229 -0.080 0.322 0.122 ;
      RECT 0.000 -0.080 0.229 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.129 1.120 1.800 1.280 ;
      RECT 1.006 1.078 1.129 1.280 ;
      RECT 0.725 1.120 1.006 1.280 ;
      RECT 0.633 1.078 0.725 1.280 ;
      RECT 0.338 1.120 0.633 1.280 ;
      RECT 0.323 1.078 0.338 1.280 ;
      RECT 0.260 1.065 0.323 1.280 ;
      RECT 0.245 1.078 0.260 1.280 ;
      RECT 0.000 1.120 0.245 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.886 0.400 0.989 0.487 ;
      RECT 0.274 0.400 0.886 0.455 ;
      RECT 0.211 0.302 0.274 0.799 ;
      RECT 0.142 0.302 0.211 0.357 ;
      RECT 0.142 0.744 0.211 0.799 ;
      RECT 0.049 0.276 0.142 0.357 ;
      RECT 0.049 0.731 0.142 0.812 ;
  END
END NAND4BX2

MACRO NAND4BX1
  CLASS CORE ;
  FOREIGN NAND4BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.240 0.573 1.265 0.933 ;
      RECT 1.200 0.201 1.240 0.933 ;
      RECT 1.175 0.201 1.200 0.627 ;
      RECT 0.746 0.879 1.200 0.933 ;
      RECT 1.154 0.201 1.175 0.306 ;
      RECT 0.837 0.201 1.154 0.256 ;
      RECT 0.741 0.201 0.837 0.282 ;
      RECT 0.681 0.737 0.746 0.933 ;
      RECT 0.650 0.737 0.681 0.839 ;
      RECT 0.597 0.763 0.650 0.839 ;
      RECT 0.363 0.763 0.597 0.818 ;
      RECT 0.267 0.737 0.363 0.818 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.252 0.439 0.311 0.494 ;
      RECT 0.187 0.439 0.252 0.600 ;
      RECT 0.162 0.492 0.187 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.466 0.439 0.497 0.494 ;
      RECT 0.443 0.439 0.466 0.623 ;
      RECT 0.401 0.439 0.443 0.636 ;
      RECT 0.348 0.555 0.401 0.636 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.567 0.555 0.743 0.665 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.075 0.498 1.089 0.579 ;
      RECT 0.950 0.498 1.075 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 -0.080 1.300 0.080 ;
      RECT 1.154 -0.080 1.249 0.122 ;
      RECT 0.151 -0.080 1.154 0.080 ;
      RECT 0.055 -0.080 0.151 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.957 1.120 1.300 1.280 ;
      RECT 0.830 1.078 0.957 1.280 ;
      RECT 0.554 1.120 0.830 1.280 ;
      RECT 0.459 1.078 0.554 1.280 ;
      RECT 0.174 1.120 0.459 1.280 ;
      RECT 0.079 1.078 0.174 1.280 ;
      RECT 0.000 1.120 0.079 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.040 0.737 1.135 0.818 ;
      RECT 0.881 0.737 1.040 0.792 ;
      RECT 0.992 0.311 1.034 0.392 ;
      RECT 0.938 0.311 0.992 0.405 ;
      RECT 0.927 0.324 0.938 0.405 ;
      RECT 0.881 0.350 0.927 0.405 ;
      RECT 0.816 0.350 0.881 0.792 ;
      RECT 0.758 0.419 0.816 0.500 ;
  END
END NAND4BX1

MACRO NAND4XL
  CLASS CORE ;
  FOREIGN NAND4XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.660 0.296 0.811 0.377 ;
      RECT 0.592 0.737 0.685 0.818 ;
      RECT 0.481 0.323 0.660 0.377 ;
      RECT 0.481 0.737 0.592 0.792 ;
      RECT 0.419 0.323 0.481 0.792 ;
      RECT 0.308 0.737 0.419 0.792 ;
      RECT 0.215 0.737 0.308 0.818 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.142 0.558 0.176 0.639 ;
      RECT 0.079 0.439 0.142 0.639 ;
      RECT 0.059 0.439 0.079 0.494 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.330 0.558 0.346 0.639 ;
      RECT 0.267 0.439 0.330 0.639 ;
      RECT 0.239 0.439 0.267 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.623 0.439 0.661 0.494 ;
      RECT 0.560 0.439 0.623 0.639 ;
      RECT 0.544 0.558 0.560 0.639 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.837 0.439 0.841 0.494 ;
      RECT 0.758 0.439 0.837 0.639 ;
      RECT 0.745 0.558 0.758 0.639 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.146 -0.080 0.900 0.080 ;
      RECT 0.053 -0.080 0.146 0.122 ;
      RECT 0.000 -0.080 0.053 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.758 1.078 0.851 1.280 ;
      RECT 0.569 1.120 0.758 1.280 ;
      RECT 0.472 1.078 0.569 1.280 ;
      RECT 0.142 1.120 0.472 1.280 ;
      RECT 0.049 1.078 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
END NAND4XL

MACRO NAND4X4
  CLASS CORE ;
  FOREIGN NAND4X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.786 0.192 2.803 0.639 ;
      RECT 2.775 0.192 2.786 0.900 ;
      RECT 2.723 0.192 2.775 0.942 ;
      RECT 2.684 0.192 2.723 0.307 ;
      RECT 2.684 0.567 2.723 0.942 ;
      RECT 2.176 0.192 2.684 0.263 ;
      RECT 2.100 0.870 2.684 0.942 ;
      RECT 2.123 0.150 2.176 0.263 ;
      RECT 2.032 0.150 2.123 0.343 ;
      RECT 0.287 0.870 2.100 0.937 ;
      RECT 0.818 0.207 2.032 0.274 ;
      RECT 0.727 0.150 0.818 0.343 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.618 0.426 2.662 0.507 ;
      RECT 2.572 0.426 2.618 0.815 ;
      RECT 2.556 0.439 2.572 0.815 ;
      RECT 1.471 0.761 2.556 0.815 ;
      RECT 1.380 0.735 1.471 0.815 ;
      RECT 0.295 0.761 1.380 0.815 ;
      RECT 0.273 0.706 0.295 0.815 ;
      RECT 0.234 0.519 0.273 0.815 ;
      RECT 0.211 0.519 0.234 0.761 ;
      RECT 0.182 0.519 0.211 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.472 0.519 2.487 0.600 ;
      RECT 2.396 0.519 2.472 0.633 ;
      RECT 2.393 0.573 2.396 0.633 ;
      RECT 2.352 0.573 2.393 0.706 ;
      RECT 2.332 0.579 2.352 0.706 ;
      RECT 1.726 0.651 2.332 0.706 ;
      RECT 1.635 0.625 1.726 0.706 ;
      RECT 1.214 0.625 1.635 0.680 ;
      RECT 1.123 0.625 1.214 0.706 ;
      RECT 0.472 0.651 1.123 0.706 ;
      RECT 0.410 0.519 0.472 0.706 ;
      RECT 0.364 0.519 0.410 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.257 0.515 2.270 0.596 ;
      RECT 2.155 0.433 2.257 0.596 ;
      RECT 1.912 0.542 2.155 0.596 ;
      RECT 1.811 0.510 1.912 0.596 ;
      RECT 1.036 0.510 1.811 0.564 ;
      RECT 0.936 0.510 1.036 0.596 ;
      RECT 0.642 0.542 0.936 0.596 ;
      RECT 0.541 0.515 0.642 0.596 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.988 0.400 2.088 0.487 ;
      RECT 0.826 0.400 1.988 0.455 ;
      RECT 0.726 0.400 0.826 0.487 ;
      RECT 0.492 0.400 0.726 0.455 ;
      RECT 0.430 0.306 0.492 0.455 ;
      RECT 0.410 0.306 0.430 0.361 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.775 -0.080 3.000 0.080 ;
      RECT 2.684 -0.080 2.775 0.122 ;
      RECT 1.471 -0.080 2.684 0.080 ;
      RECT 1.380 -0.080 1.471 0.122 ;
      RECT 0.166 -0.080 1.380 0.080 ;
      RECT 0.075 -0.080 0.166 0.122 ;
      RECT 0.000 -0.080 0.075 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.753 1.120 3.000 1.280 ;
      RECT 2.662 1.078 2.753 1.280 ;
      RECT 2.373 1.120 2.662 1.280 ;
      RECT 2.282 1.078 2.373 1.280 ;
      RECT 2.007 1.120 2.282 1.280 ;
      RECT 1.886 1.078 2.007 1.280 ;
      RECT 0.964 1.120 1.886 1.280 ;
      RECT 0.844 1.078 0.964 1.280 ;
      RECT 0.568 1.120 0.844 1.280 ;
      RECT 0.477 1.078 0.568 1.280 ;
      RECT 0.189 1.120 0.477 1.280 ;
      RECT 0.098 1.078 0.189 1.280 ;
      RECT 0.000 1.120 0.098 1.280 ;
     END
  END VDD
END NAND4X4

MACRO NAND4X2
  CLASS CORE ;
  FOREIGN NAND4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 0.195 1.542 0.633 ;
      RECT 1.467 0.195 1.541 0.973 ;
      RECT 1.460 0.195 1.467 0.306 ;
      RECT 1.460 0.564 1.467 0.973 ;
      RECT 0.797 0.195 1.460 0.262 ;
      RECT 0.854 0.901 1.460 0.973 ;
      RECT 0.773 0.870 0.854 0.973 ;
      RECT 0.706 0.150 0.797 0.343 ;
      RECT 0.256 0.870 0.773 0.942 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.162 0.761 1.254 0.842 ;
      RECT 0.298 0.761 1.162 0.815 ;
      RECT 0.241 0.706 0.298 0.815 ;
      RECT 0.236 0.519 0.241 0.815 ;
      RECT 0.179 0.519 0.236 0.761 ;
      RECT 0.149 0.519 0.179 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.187 0.519 1.193 0.600 ;
      RECT 1.164 0.519 1.187 0.627 ;
      RECT 1.102 0.519 1.164 0.706 ;
      RECT 0.442 0.651 1.102 0.706 ;
      RECT 0.380 0.519 0.442 0.706 ;
      RECT 0.333 0.519 0.380 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.916 0.439 1.017 0.596 ;
      RECT 0.613 0.542 0.916 0.596 ;
      RECT 0.512 0.515 0.613 0.596 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.698 0.401 0.799 0.487 ;
      RECT 0.496 0.401 0.698 0.456 ;
      RECT 0.434 0.306 0.496 0.456 ;
      RECT 0.413 0.306 0.434 0.361 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.455 -0.080 1.600 0.080 ;
      RECT 1.363 -0.080 1.455 0.122 ;
      RECT 0.140 -0.080 1.363 0.080 ;
      RECT 0.048 -0.080 0.140 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.937 1.120 1.600 1.280 ;
      RECT 0.816 1.078 0.937 1.280 ;
      RECT 0.539 1.120 0.816 1.280 ;
      RECT 0.447 1.078 0.539 1.280 ;
      RECT 0.156 1.120 0.447 1.280 ;
      RECT 0.065 1.078 0.156 1.280 ;
      RECT 0.000 1.120 0.065 1.280 ;
     END
  END VDD
END NAND4X2

MACRO NAND4X1
  CLASS CORE ;
  FOREIGN NAND4X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.817 0.308 0.865 0.792 ;
      RECT 0.802 0.170 0.817 0.792 ;
      RECT 0.724 0.170 0.802 0.363 ;
      RECT 0.758 0.706 0.802 0.792 ;
      RECT 0.682 0.737 0.758 0.792 ;
      RECT 0.589 0.737 0.682 0.818 ;
      RECT 0.311 0.737 0.589 0.792 ;
      RECT 0.218 0.737 0.311 0.818 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.142 0.555 0.210 0.636 ;
      RECT 0.079 0.439 0.142 0.636 ;
      RECT 0.059 0.439 0.079 0.494 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.335 0.555 0.405 0.636 ;
      RECT 0.273 0.439 0.335 0.636 ;
      RECT 0.239 0.439 0.273 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.521 0.573 0.682 0.662 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.645 0.419 0.738 0.500 ;
      RECT 0.419 0.439 0.645 0.494 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.146 -0.080 0.900 0.080 ;
      RECT 0.053 -0.080 0.146 0.247 ;
      RECT 0.000 -0.080 0.053 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.758 1.078 0.851 1.280 ;
      RECT 0.567 1.120 0.758 1.280 ;
      RECT 0.475 1.078 0.567 1.280 ;
      RECT 0.142 1.120 0.475 1.280 ;
      RECT 0.049 1.078 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
END NAND4X1

MACRO NAND3BXL
  CLASS CORE ;
  FOREIGN NAND3BXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.158 0.862 1.042 ;
      RECT 0.742 0.158 0.799 0.213 ;
      RECT 0.779 0.700 0.799 1.042 ;
      RECT 0.758 0.700 0.779 0.854 ;
      RECT 0.753 0.987 0.779 1.042 ;
      RECT 0.502 0.799 0.758 0.854 ;
      RECT 0.409 0.786 0.502 0.867 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.331 0.607 0.393 0.719 ;
      RECT 0.330 0.607 0.331 0.767 ;
      RECT 0.218 0.664 0.330 0.767 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.379 0.581 0.500 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.367 0.142 0.500 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.322 -0.080 0.900 0.080 ;
      RECT 0.229 -0.080 0.322 0.122 ;
      RECT 0.000 -0.080 0.229 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.655 1.120 0.900 1.280 ;
      RECT 0.562 1.078 0.655 1.280 ;
      RECT 0.322 1.120 0.562 1.280 ;
      RECT 0.229 1.078 0.322 1.280 ;
      RECT 0.000 1.120 0.229 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.672 0.268 0.735 0.607 ;
      RECT 0.267 0.268 0.672 0.323 ;
      RECT 0.205 0.257 0.267 0.610 ;
      RECT 0.049 0.257 0.205 0.312 ;
      RECT 0.127 0.555 0.205 0.610 ;
      RECT 0.127 0.764 0.142 0.845 ;
      RECT 0.064 0.555 0.127 0.845 ;
      RECT 0.049 0.764 0.064 0.845 ;
  END
END NAND3BXL

MACRO NAND3BX4
  CLASS CORE ;
  FOREIGN NAND3BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.887 0.199 1.950 0.755 ;
      RECT 1.846 0.199 1.887 0.307 ;
      RECT 1.780 0.700 1.887 0.755 ;
      RECT 0.882 0.199 1.846 0.254 ;
      RECT 1.723 0.700 1.780 1.033 ;
      RECT 1.675 0.688 1.723 1.033 ;
      RECT 1.577 0.688 1.675 0.810 ;
      RECT 0.977 0.755 1.577 0.810 ;
      RECT 0.883 0.742 0.977 0.823 ;
      RECT 0.850 0.742 0.883 0.810 ;
      RECT 0.788 0.167 0.882 0.254 ;
      RECT 0.585 0.755 0.850 0.810 ;
      RECT 0.492 0.742 0.585 0.823 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.234 0.915 1.328 0.996 ;
      RECT 0.397 0.929 1.234 0.983 ;
      RECT 0.397 0.439 0.486 0.500 ;
      RECT 0.333 0.439 0.397 0.983 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.489 0.507 1.583 0.607 ;
      RECT 1.234 0.507 1.489 0.562 ;
      RECT 1.132 0.507 1.234 0.633 ;
      RECT 1.039 0.494 1.132 0.633 ;
      RECT 1.032 0.567 1.039 0.633 ;
      RECT 0.661 0.579 1.032 0.633 ;
      RECT 0.567 0.577 0.661 0.658 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.047 0.411 0.140 0.563 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.405 -0.080 2.000 0.080 ;
      RECT 1.311 -0.080 1.405 0.122 ;
      RECT 0.358 -0.080 1.311 0.080 ;
      RECT 0.264 -0.080 0.358 0.122 ;
      RECT 0.000 -0.080 0.264 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.906 1.120 2.000 1.280 ;
      RECT 1.843 0.905 1.906 1.280 ;
      RECT 1.528 1.120 1.843 1.280 ;
      RECT 1.434 0.905 1.528 1.280 ;
      RECT 1.164 1.120 1.434 1.280 ;
      RECT 1.070 1.078 1.164 1.280 ;
      RECT 0.781 1.120 1.070 1.280 ;
      RECT 0.687 1.078 0.781 1.280 ;
      RECT 0.362 1.120 0.687 1.280 ;
      RECT 0.269 1.078 0.362 1.280 ;
      RECT 0.000 1.120 0.269 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.775 0.440 1.822 0.555 ;
      RECT 1.759 0.315 1.775 0.555 ;
      RECT 1.712 0.315 1.759 0.495 ;
      RECT 0.848 0.315 1.712 0.370 ;
      RECT 0.755 0.315 0.848 0.496 ;
      RECT 0.270 0.315 0.755 0.370 ;
      RECT 0.207 0.250 0.270 0.745 ;
      RECT 0.143 0.250 0.207 0.305 ;
      RECT 0.143 0.690 0.207 0.745 ;
      RECT 0.050 0.224 0.143 0.305 ;
      RECT 0.050 0.690 0.143 0.771 ;
  END
END NAND3BX4

MACRO NAND3BX2
  CLASS CORE ;
  FOREIGN NAND3BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.651 0.689 0.741 0.770 ;
      RECT 0.567 0.164 0.658 0.245 ;
      RECT 0.643 0.689 0.651 0.767 ;
      RECT 0.407 0.700 0.643 0.767 ;
      RECT 0.294 0.177 0.567 0.232 ;
      RECT 0.373 0.689 0.407 0.767 ;
      RECT 0.294 0.689 0.373 0.770 ;
      RECT 0.282 0.177 0.294 0.770 ;
      RECT 0.233 0.177 0.282 0.767 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.033 0.462 1.047 0.543 ;
      RECT 0.972 0.462 1.033 0.881 ;
      RECT 0.957 0.462 0.972 0.543 ;
      RECT 0.172 0.826 0.972 0.881 ;
      RECT 0.111 0.439 0.172 0.881 ;
      RECT 0.082 0.439 0.111 0.573 ;
      RECT 0.057 0.439 0.082 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.838 0.507 0.870 0.588 ;
      RECT 0.737 0.433 0.838 0.604 ;
      RECT 0.445 0.549 0.737 0.604 ;
      RECT 0.355 0.514 0.445 0.604 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.358 0.467 1.363 0.594 ;
      RECT 1.267 0.433 1.358 0.594 ;
      RECT 1.262 0.467 1.267 0.594 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.161 -0.080 1.400 0.080 ;
      RECT 1.145 -0.080 1.161 0.122 ;
      RECT 1.055 -0.080 1.145 0.247 ;
      RECT 0.154 -0.080 1.055 0.080 ;
      RECT 0.064 -0.080 0.154 0.247 ;
      RECT 0.000 -0.080 0.064 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.148 1.120 1.400 1.280 ;
      RECT 1.058 0.952 1.148 1.280 ;
      RECT 0.561 1.120 1.058 1.280 ;
      RECT 0.471 0.952 0.561 1.280 ;
      RECT 0.192 1.120 0.471 1.280 ;
      RECT 0.102 0.952 0.192 1.280 ;
      RECT 0.000 1.120 0.102 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.262 0.279 1.352 0.379 ;
      RECT 1.262 0.702 1.352 0.783 ;
      RECT 1.201 0.324 1.262 0.379 ;
      RECT 1.201 0.702 1.262 0.757 ;
      RECT 1.140 0.324 1.201 0.757 ;
      RECT 0.658 0.324 1.140 0.379 ;
      RECT 0.597 0.324 0.658 0.490 ;
      RECT 0.567 0.410 0.597 0.490 ;
  END
END NAND3BX2

MACRO NAND3BX1
  CLASS CORE ;
  FOREIGN NAND3BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.158 0.862 1.042 ;
      RECT 0.742 0.158 0.799 0.213 ;
      RECT 0.779 0.833 0.799 1.042 ;
      RECT 0.502 0.833 0.779 0.888 ;
      RECT 0.753 0.987 0.779 1.042 ;
      RECT 0.409 0.833 0.502 0.914 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.330 0.593 0.393 0.761 ;
      RECT 0.239 0.665 0.330 0.761 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.414 0.567 0.500 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.367 0.142 0.500 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.305 -0.080 0.900 0.080 ;
      RECT 0.213 -0.080 0.305 0.122 ;
      RECT 0.000 -0.080 0.213 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.655 1.120 0.900 1.280 ;
      RECT 0.562 1.078 0.655 1.280 ;
      RECT 0.322 1.120 0.562 1.280 ;
      RECT 0.229 1.078 0.322 1.280 ;
      RECT 0.000 1.120 0.229 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.672 0.268 0.735 0.605 ;
      RECT 0.267 0.268 0.672 0.323 ;
      RECT 0.205 0.257 0.267 0.610 ;
      RECT 0.049 0.257 0.205 0.312 ;
      RECT 0.127 0.555 0.205 0.610 ;
      RECT 0.127 0.854 0.142 0.935 ;
      RECT 0.064 0.555 0.127 0.935 ;
      RECT 0.049 0.854 0.064 0.935 ;
  END
END NAND3BX1

MACRO NAND3XL
  CLASS CORE ;
  FOREIGN NAND3XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.591 0.251 0.652 0.782 ;
      RECT 0.562 0.251 0.591 0.332 ;
      RECT 0.562 0.681 0.591 0.782 ;
      RECT 0.278 0.727 0.562 0.782 ;
      RECT 0.188 0.714 0.278 0.795 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.487 0.138 0.633 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.433 0.349 0.617 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.500 0.536 0.529 0.617 ;
      RECT 0.439 0.306 0.500 0.617 ;
      RECT 0.407 0.306 0.439 0.361 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.138 -0.080 0.700 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.456 1.120 0.700 1.280 ;
      RECT 0.119 1.078 0.456 1.280 ;
      RECT 0.000 1.120 0.119 1.280 ;
     END
  END VDD
END NAND3XL

MACRO NAND3X4
  CLASS CORE ;
  FOREIGN NAND3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.707 0.158 1.713 0.351 ;
      RECT 1.645 0.158 1.707 0.744 ;
      RECT 1.620 0.158 1.645 0.351 ;
      RECT 1.510 0.689 1.645 0.744 ;
      RECT 1.560 0.158 1.620 0.248 ;
      RECT 0.676 0.193 1.560 0.248 ;
      RECT 1.417 0.689 1.510 0.770 ;
      RECT 0.316 0.689 0.770 0.770 ;
      RECT 0.322 0.167 0.676 0.248 ;
      RECT 0.316 0.167 0.322 0.500 ;
      RECT 0.224 0.167 0.316 0.770 ;
      RECT 0.218 0.167 0.224 0.500 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.098 0.527 1.113 0.608 ;
      RECT 1.035 0.527 1.098 0.880 ;
      RECT 1.020 0.527 1.035 0.608 ;
      RECT 0.155 0.825 1.035 0.880 ;
      RECT 0.093 0.439 0.155 0.880 ;
      RECT 0.059 0.439 0.093 0.573 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.365 0.494 1.395 0.590 ;
      RECT 1.302 0.418 1.365 0.590 ;
      RECT 0.927 0.418 1.302 0.473 ;
      RECT 0.835 0.417 0.927 0.498 ;
      RECT 0.821 0.418 0.835 0.498 ;
      RECT 0.758 0.418 0.821 0.601 ;
      RECT 0.477 0.546 0.758 0.601 ;
      RECT 0.385 0.514 0.477 0.601 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.546 0.426 1.579 0.590 ;
      RECT 1.486 0.302 1.546 0.590 ;
      RECT 1.484 0.302 1.486 0.499 ;
      RECT 0.676 0.302 1.484 0.357 ;
      RECT 0.614 0.302 0.676 0.492 ;
      RECT 0.584 0.411 0.614 0.492 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.195 -0.080 1.800 0.080 ;
      RECT 1.102 -0.080 1.195 0.122 ;
      RECT 0.155 -0.080 1.102 0.080 ;
      RECT 0.063 -0.080 0.155 0.247 ;
      RECT 0.000 -0.080 0.063 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.695 1.120 1.800 1.280 ;
      RECT 1.602 0.952 1.695 1.280 ;
      RECT 1.324 1.120 1.602 1.280 ;
      RECT 1.231 0.952 1.324 1.280 ;
      RECT 0.956 1.120 1.231 1.280 ;
      RECT 0.863 0.952 0.956 1.280 ;
      RECT 0.577 1.120 0.863 1.280 ;
      RECT 0.484 0.952 0.577 1.280 ;
      RECT 0.198 1.120 0.484 1.280 ;
      RECT 0.105 0.952 0.198 1.280 ;
      RECT 0.000 1.120 0.105 1.280 ;
     END
  END VDD
END NAND3X4

MACRO NAND3X2
  CLASS CORE ;
  FOREIGN NAND3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.691 0.689 0.786 0.770 ;
      RECT 0.602 0.164 0.698 0.245 ;
      RECT 0.682 0.689 0.691 0.761 ;
      RECT 0.518 0.706 0.682 0.761 ;
      RECT 0.312 0.190 0.602 0.245 ;
      RECT 0.432 0.700 0.518 0.770 ;
      RECT 0.312 0.689 0.432 0.770 ;
      RECT 0.300 0.190 0.312 0.770 ;
      RECT 0.248 0.190 0.300 0.761 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.096 0.573 1.111 0.706 ;
      RECT 1.031 0.573 1.096 0.881 ;
      RECT 1.016 0.573 1.031 0.706 ;
      RECT 0.183 0.826 1.031 0.881 ;
      RECT 0.167 0.460 0.183 0.881 ;
      RECT 0.118 0.439 0.167 0.881 ;
      RECT 0.087 0.439 0.118 0.573 ;
      RECT 0.060 0.439 0.087 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.907 0.493 0.923 0.588 ;
      RECT 0.868 0.433 0.907 0.588 ;
      RECT 0.782 0.433 0.868 0.604 ;
      RECT 0.473 0.549 0.782 0.604 ;
      RECT 0.377 0.514 0.473 0.604 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.602 0.300 0.698 0.490 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.232 -0.080 1.300 0.080 ;
      RECT 1.137 -0.080 1.232 0.122 ;
      RECT 0.163 -0.080 1.137 0.080 ;
      RECT 0.068 -0.080 0.163 0.122 ;
      RECT 0.000 -0.080 0.068 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.595 1.120 1.300 1.280 ;
      RECT 0.499 0.952 0.595 1.280 ;
      RECT 0.204 1.120 0.499 1.280 ;
      RECT 0.108 0.952 0.204 1.280 ;
      RECT 0.000 1.120 0.108 1.280 ;
     END
  END VDD
END NAND3X2

MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 0.695 0.655 0.812 ;
      RECT 0.591 0.167 0.652 0.812 ;
      RECT 0.562 0.167 0.591 0.307 ;
      RECT 0.581 0.695 0.591 0.812 ;
      RECT 0.562 0.731 0.581 0.812 ;
      RECT 0.293 0.744 0.562 0.799 ;
      RECT 0.203 0.731 0.293 0.812 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.050 0.425 0.141 0.590 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.544 0.349 0.676 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.500 0.501 0.529 0.582 ;
      RECT 0.439 0.306 0.500 0.582 ;
      RECT 0.407 0.306 0.439 0.361 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.154 -0.080 0.700 0.080 ;
      RECT 0.064 -0.080 0.154 0.122 ;
      RECT 0.000 -0.080 0.064 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.483 1.120 0.700 1.280 ;
      RECT 0.048 1.078 0.483 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
END NAND3X1

MACRO NAND2BXL
  CLASS CORE ;
  FOREIGN NAND2BXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.647 0.306 0.662 0.845 ;
      RECT 0.601 0.245 0.647 0.845 ;
      RECT 0.557 0.245 0.601 0.361 ;
      RECT 0.488 0.790 0.601 0.845 ;
      RECT 0.407 0.306 0.557 0.361 ;
      RECT 0.398 0.777 0.488 0.858 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.377 0.460 0.391 0.544 ;
      RECT 0.232 0.439 0.377 0.544 ;
      RECT 0.212 0.460 0.232 0.544 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.056 0.901 0.196 1.033 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.636 1.120 0.700 1.280 ;
      RECT 0.377 1.078 0.636 1.280 ;
      RECT 0.000 1.120 0.377 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.476 0.613 0.537 0.723 ;
      RECT 0.138 0.668 0.476 0.723 ;
      RECT 0.123 0.274 0.138 0.355 ;
      RECT 0.123 0.668 0.138 0.821 ;
      RECT 0.062 0.274 0.123 0.821 ;
      RECT 0.048 0.274 0.062 0.355 ;
      RECT 0.048 0.740 0.062 0.821 ;
  END
END NAND2BXL

MACRO NAND2BX4
  CLASS CORE ;
  FOREIGN NAND2BX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.358 0.245 1.363 0.633 ;
      RECT 1.267 0.245 1.358 0.798 ;
      RECT 1.262 0.245 1.267 0.633 ;
      RECT 0.396 0.717 1.267 0.798 ;
      RECT 0.673 0.327 1.262 0.399 ;
      RECT 0.583 0.283 0.673 0.399 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.818 0.568 0.985 0.662 ;
      RECT 0.480 0.607 0.818 0.662 ;
      RECT 0.424 0.573 0.480 0.662 ;
      RECT 0.334 0.568 0.424 0.662 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.045 0.481 0.135 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.013 -0.080 1.400 0.080 ;
      RECT 0.923 -0.080 1.013 0.254 ;
      RECT 0.339 -0.080 0.923 0.080 ;
      RECT 0.249 -0.080 0.339 0.122 ;
      RECT 0.000 -0.080 0.249 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 1.120 1.400 1.280 ;
      RECT 1.246 0.871 1.336 1.280 ;
      RECT 0.996 1.120 1.246 1.280 ;
      RECT 0.905 0.871 0.996 1.280 ;
      RECT 0.656 1.120 0.905 1.280 ;
      RECT 0.566 0.871 0.656 1.280 ;
      RECT 0.317 1.120 0.566 1.280 ;
      RECT 0.227 0.883 0.317 1.280 ;
      RECT 0.000 1.120 0.227 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.140 0.457 1.201 0.649 ;
      RECT 0.671 0.457 1.140 0.512 ;
      RECT 0.581 0.457 0.671 0.552 ;
      RECT 0.260 0.457 0.581 0.512 ;
      RECT 0.199 0.305 0.260 0.771 ;
      RECT 0.138 0.305 0.199 0.360 ;
      RECT 0.138 0.717 0.199 0.771 ;
      RECT 0.048 0.279 0.138 0.360 ;
      RECT 0.048 0.717 0.138 0.798 ;
  END
END NAND2BX4

MACRO NAND2BX2
  CLASS CORE ;
  FOREIGN NAND2BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.003 0.402 1.067 0.770 ;
      RECT 0.878 0.402 1.003 0.457 ;
      RECT 0.894 0.700 1.003 0.770 ;
      RECT 0.800 0.690 0.894 0.771 ;
      RECT 0.876 0.361 0.878 0.457 ;
      RECT 0.812 0.317 0.876 0.457 ;
      RECT 0.694 0.317 0.812 0.371 ;
      RECT 0.772 0.700 0.800 0.770 ;
      RECT 0.610 0.715 0.772 0.770 ;
      RECT 0.600 0.290 0.694 0.371 ;
      RECT 0.539 0.702 0.610 0.770 ;
      RECT 0.444 0.702 0.539 0.783 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.853 0.549 0.939 0.636 ;
      RECT 0.467 0.573 0.853 0.627 ;
      RECT 0.372 0.560 0.467 0.640 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.047 0.452 0.142 0.627 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 -0.080 1.100 0.080 ;
      RECT 0.956 -0.080 1.050 0.278 ;
      RECT 0.328 -0.080 0.956 0.080 ;
      RECT 0.233 -0.080 0.328 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 1.120 1.100 1.280 ;
      RECT 0.353 1.078 1.050 1.280 ;
      RECT 0.000 1.120 0.353 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.639 0.433 0.733 0.514 ;
      RECT 0.272 0.446 0.639 0.501 ;
      RECT 0.208 0.311 0.272 0.757 ;
      RECT 0.144 0.311 0.208 0.368 ;
      RECT 0.144 0.702 0.208 0.757 ;
      RECT 0.050 0.279 0.144 0.368 ;
      RECT 0.050 0.702 0.144 0.783 ;
      RECT 0.049 0.292 0.050 0.368 ;
  END
END NAND2BX2

MACRO NAND2BX1
  CLASS CORE ;
  FOREIGN NAND2BX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.586 0.289 0.647 0.808 ;
      RECT 0.557 0.289 0.586 0.370 ;
      RECT 0.398 0.754 0.586 0.808 ;
      RECT 0.467 0.300 0.557 0.367 ;
      RECT 0.407 0.306 0.467 0.361 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.377 0.461 0.391 0.545 ;
      RECT 0.232 0.439 0.377 0.545 ;
      RECT 0.212 0.461 0.232 0.545 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.056 0.901 0.196 1.033 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.636 1.120 0.700 1.280 ;
      RECT 0.377 1.078 0.636 1.280 ;
      RECT 0.000 1.120 0.377 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.463 0.605 0.524 0.694 ;
      RECT 0.123 0.605 0.463 0.660 ;
      RECT 0.123 0.274 0.138 0.355 ;
      RECT 0.123 0.740 0.138 0.821 ;
      RECT 0.062 0.274 0.123 0.821 ;
      RECT 0.048 0.274 0.062 0.355 ;
      RECT 0.048 0.740 0.062 0.821 ;
  END
END NAND2BX1

MACRO NAND2XL
  CLASS CORE ;
  FOREIGN NAND2XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.545 0.294 0.552 0.770 ;
      RECT 0.535 0.281 0.545 0.770 ;
      RECT 0.482 0.281 0.535 0.798 ;
      RECT 0.442 0.281 0.482 0.362 ;
      RECT 0.452 0.695 0.482 0.798 ;
      RECT 0.355 0.743 0.452 0.798 ;
      RECT 0.252 0.743 0.355 0.824 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.500 0.158 0.645 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.379 0.494 0.412 0.624 ;
      RECT 0.309 0.439 0.379 0.624 ;
      RECT 0.265 0.439 0.309 0.494 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 -0.080 0.600 0.080 ;
      RECT 0.055 -0.080 0.158 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.321 1.120 0.600 1.280 ;
      RECT 0.148 1.078 0.321 1.280 ;
      RECT 0.000 1.120 0.148 1.280 ;
     END
  END VDD
END NAND2XL

MACRO NAND2X4
  CLASS CORE ;
  FOREIGN NAND2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 0.245 1.261 0.633 ;
      RECT 1.154 0.245 1.249 0.798 ;
      RECT 0.529 0.307 1.154 0.379 ;
      RECT 0.231 0.717 1.154 0.798 ;
      RECT 0.433 0.283 0.529 0.379 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.844 0.576 0.860 0.657 ;
      RECT 0.764 0.576 0.844 0.662 ;
      RECT 0.311 0.607 0.764 0.662 ;
      RECT 0.184 0.573 0.311 0.662 ;
      RECT 0.169 0.573 0.184 0.654 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.024 0.467 1.089 0.652 ;
      RECT 0.968 0.467 1.024 0.573 ;
      RECT 0.695 0.467 0.968 0.521 ;
      RECT 0.605 0.439 0.695 0.521 ;
      RECT 0.526 0.467 0.605 0.521 ;
      RECT 0.446 0.467 0.526 0.552 ;
      RECT 0.431 0.471 0.446 0.552 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.889 -0.080 1.300 0.080 ;
      RECT 0.794 -0.080 0.889 0.237 ;
      RECT 0.174 -0.080 0.794 0.080 ;
      RECT 0.079 -0.080 0.174 0.122 ;
      RECT 0.000 -0.080 0.079 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.227 1.120 1.300 1.280 ;
      RECT 1.131 0.871 1.227 1.280 ;
      RECT 0.867 1.120 1.131 1.280 ;
      RECT 0.771 0.871 0.867 1.280 ;
      RECT 0.506 1.120 0.771 1.280 ;
      RECT 0.411 0.871 0.506 1.280 ;
      RECT 0.146 1.120 0.411 1.280 ;
      RECT 0.051 0.871 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
END NAND2X4

MACRO NAND2X2
  CLASS CORE ;
  FOREIGN NAND2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.795 0.402 0.858 0.770 ;
      RECT 0.680 0.402 0.795 0.457 ;
      RECT 0.779 0.704 0.795 0.770 ;
      RECT 0.251 0.704 0.779 0.758 ;
      RECT 0.618 0.249 0.680 0.457 ;
      RECT 0.599 0.249 0.618 0.306 ;
      RECT 0.502 0.249 0.599 0.304 ;
      RECT 0.409 0.223 0.502 0.304 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.668 0.558 0.731 0.645 ;
      RECT 0.301 0.577 0.668 0.632 ;
      RECT 0.200 0.573 0.301 0.632 ;
      RECT 0.185 0.573 0.200 0.627 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.400 0.551 0.520 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.289 ;
      RECT 0.142 -0.080 0.758 0.080 ;
      RECT 0.049 -0.080 0.142 0.122 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.210 1.078 0.851 1.280 ;
      RECT 0.000 1.120 0.210 1.280 ;
     END
  END VDD
END NAND2X2

MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.545 0.300 0.564 0.743 ;
      RECT 0.494 0.282 0.545 0.743 ;
      RECT 0.442 0.282 0.494 0.367 ;
      RECT 0.352 0.688 0.494 0.743 ;
      RECT 0.248 0.688 0.352 0.769 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.438 0.158 0.598 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.242 0.530 0.421 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 -0.080 0.600 0.080 ;
      RECT 0.055 -0.080 0.158 0.328 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.359 1.120 0.600 1.280 ;
      RECT 0.055 1.078 0.359 1.280 ;
      RECT 0.000 1.120 0.055 1.280 ;
     END
  END VDD
END NAND2X1

MACRO MXI4X4
  CLASS CORE ;
  FOREIGN MXI4X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.101 0.235 4.187 0.904 ;
      RECT 4.085 0.183 4.101 1.015 ;
      RECT 4.011 0.183 4.085 0.376 ;
      RECT 4.011 0.711 4.085 1.015 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.205 0.550 3.355 0.640 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.093 0.433 1.205 0.567 ;
     END
  END S0

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.500 0.433 1.547 0.500 ;
      RECT 1.399 0.433 1.500 0.546 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.291 0.300 2.412 0.367 ;
      RECT 2.231 0.300 2.291 0.561 ;
      RECT 2.229 0.306 2.231 0.561 ;
      RECT 2.203 0.474 2.229 0.561 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.019 0.469 1.025 0.546 ;
      RECT 0.917 0.302 1.019 0.546 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.526 0.208 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.304 -0.080 4.400 0.080 ;
      RECT 4.213 -0.080 4.304 0.122 ;
      RECT 3.899 -0.080 4.213 0.080 ;
      RECT 3.808 -0.080 3.899 0.122 ;
      RECT 3.509 -0.080 3.808 0.080 ;
      RECT 3.419 -0.080 3.509 0.122 ;
      RECT 2.359 -0.080 3.419 0.080 ;
      RECT 2.268 -0.080 2.359 0.217 ;
      RECT 1.465 -0.080 2.268 0.080 ;
      RECT 1.375 -0.080 1.465 0.230 ;
      RECT 1.059 -0.080 1.375 0.080 ;
      RECT 0.968 -0.080 1.059 0.220 ;
      RECT 0.152 -0.080 0.968 0.080 ;
      RECT 0.061 -0.080 0.152 0.289 ;
      RECT 0.000 -0.080 0.061 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.304 1.120 4.400 1.280 ;
      RECT 4.213 1.078 4.304 1.280 ;
      RECT 3.899 1.120 4.213 1.280 ;
      RECT 3.808 1.078 3.899 1.280 ;
      RECT 3.461 1.120 3.808 1.280 ;
      RECT 3.371 1.078 3.461 1.280 ;
      RECT 2.359 1.120 3.371 1.280 ;
      RECT 2.268 1.078 2.359 1.280 ;
      RECT 1.463 1.120 2.268 1.280 ;
      RECT 1.372 0.998 1.463 1.280 ;
      RECT 1.059 1.120 1.372 1.280 ;
      RECT 0.968 0.998 1.059 1.280 ;
      RECT 0.152 1.120 0.968 1.280 ;
      RECT 0.061 0.866 0.152 1.280 ;
      RECT 0.000 1.120 0.061 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.944 0.496 3.973 0.577 ;
      RECT 3.883 0.198 3.944 0.577 ;
      RECT 3.315 0.198 3.883 0.252 ;
      RECT 3.735 0.540 3.796 1.008 ;
      RECT 3.696 0.540 3.735 0.595 ;
      RECT 1.655 0.954 3.735 1.008 ;
      RECT 3.524 0.313 3.712 0.368 ;
      RECT 3.605 0.514 3.696 0.595 ;
      RECT 3.524 0.705 3.669 0.898 ;
      RECT 3.463 0.313 3.524 0.898 ;
      RECT 2.988 0.843 3.463 0.898 ;
      RECT 3.253 0.163 3.315 0.252 ;
      RECT 3.144 0.338 3.257 0.393 ;
      RECT 2.769 0.163 3.253 0.218 ;
      RECT 3.144 0.733 3.248 0.788 ;
      RECT 3.083 0.338 3.144 0.788 ;
      RECT 2.936 0.796 2.988 0.898 ;
      RECT 2.936 0.365 2.949 0.452 ;
      RECT 2.875 0.365 2.936 0.898 ;
      RECT 2.755 0.796 2.781 0.877 ;
      RECT 2.755 0.163 2.769 0.317 ;
      RECT 2.708 0.163 2.755 0.877 ;
      RECT 2.693 0.236 2.708 0.877 ;
      RECT 2.679 0.236 2.693 0.317 ;
      RECT 2.528 0.177 2.589 0.876 ;
      RECT 2.465 0.177 2.528 0.232 ;
      RECT 2.400 0.495 2.461 0.898 ;
      RECT 1.943 0.843 2.400 0.898 ;
      RECT 2.008 0.339 2.069 0.735 ;
      RECT 1.881 0.176 1.943 0.898 ;
      RECT 1.768 0.176 1.881 0.231 ;
      RECT 1.759 0.843 1.881 0.898 ;
      RECT 1.756 0.324 1.817 0.765 ;
      RECT 1.580 0.324 1.756 0.379 ;
      RECT 1.556 0.711 1.756 0.765 ;
      RECT 1.595 0.552 1.695 0.656 ;
      RECT 1.593 0.874 1.655 1.008 ;
      RECT 1.328 0.601 1.595 0.656 ;
      RECT 0.599 0.874 1.593 0.929 ;
      RECT 1.267 0.296 1.328 0.744 ;
      RECT 1.176 0.296 1.267 0.377 ;
      RECT 1.019 0.689 1.267 0.744 ;
      RECT 0.957 0.601 1.019 0.744 ;
      RECT 0.824 0.601 0.957 0.656 ;
      RECT 0.701 0.711 0.861 0.765 ;
      RECT 0.784 0.343 0.856 0.433 ;
      RECT 0.763 0.526 0.824 0.656 ;
      RECT 0.701 0.379 0.784 0.433 ;
      RECT 0.640 0.379 0.701 0.765 ;
      RECT 0.569 0.223 0.653 0.304 ;
      RECT 0.569 0.848 0.599 0.929 ;
      RECT 0.508 0.223 0.569 0.929 ;
      RECT 0.331 0.226 0.387 0.426 ;
      RECT 0.269 0.226 0.331 0.736 ;
  END
END MXI4X4

MACRO MXI4X2
  CLASS CORE ;
  FOREIGN MXI4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.087 0.183 4.148 1.007 ;
      RECT 4.052 0.183 4.087 0.376 ;
      RECT 4.082 0.627 4.087 1.007 ;
      RECT 4.049 0.665 4.082 1.007 ;
      RECT 3.887 0.665 4.049 0.767 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.187 0.433 3.371 0.524 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.053 0.433 1.188 0.567 ;
     END
  END S0

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.437 0.302 1.548 0.533 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.292 0.300 2.413 0.367 ;
      RECT 2.233 0.300 2.292 0.561 ;
      RECT 2.231 0.306 2.233 0.561 ;
      RECT 2.205 0.474 2.231 0.561 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.969 0.306 0.993 0.361 ;
      RECT 0.908 0.306 0.969 0.527 ;
      RECT 0.862 0.450 0.908 0.527 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.526 0.209 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.924 -0.080 4.200 0.080 ;
      RECT 3.834 -0.080 3.924 0.122 ;
      RECT 3.468 -0.080 3.834 0.080 ;
      RECT 3.378 -0.080 3.468 0.122 ;
      RECT 2.360 -0.080 3.378 0.080 ;
      RECT 2.270 -0.080 2.360 0.217 ;
      RECT 1.522 -0.080 2.270 0.080 ;
      RECT 1.432 -0.080 1.522 0.217 ;
      RECT 1.042 -0.080 1.432 0.080 ;
      RECT 0.952 -0.080 1.042 0.220 ;
      RECT 0.151 -0.080 0.952 0.080 ;
      RECT 0.061 -0.080 0.151 0.329 ;
      RECT 0.000 -0.080 0.061 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.900 1.120 4.200 1.280 ;
      RECT 3.810 1.078 3.900 1.280 ;
      RECT 3.434 1.120 3.810 1.280 ;
      RECT 3.344 1.078 3.434 1.280 ;
      RECT 2.360 1.120 3.344 1.280 ;
      RECT 2.270 1.078 2.360 1.280 ;
      RECT 1.469 1.120 2.270 1.280 ;
      RECT 1.379 0.954 1.469 1.280 ;
      RECT 1.042 1.120 1.379 1.280 ;
      RECT 0.952 0.954 1.042 1.280 ;
      RECT 0.151 1.120 0.952 1.280 ;
      RECT 0.061 0.745 0.151 1.280 ;
      RECT 0.000 1.120 0.061 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.975 0.496 4.004 0.577 ;
      RECT 3.914 0.198 3.975 0.577 ;
      RECT 3.310 0.198 3.914 0.252 ;
      RECT 3.716 0.542 3.777 1.008 ;
      RECT 3.509 0.313 3.717 0.368 ;
      RECT 3.680 0.542 3.716 0.596 ;
      RECT 1.645 0.954 3.716 1.008 ;
      RECT 3.605 0.514 3.680 0.596 ;
      RECT 3.509 0.761 3.639 0.854 ;
      RECT 3.590 0.514 3.605 0.595 ;
      RECT 3.448 0.313 3.509 0.854 ;
      RECT 2.986 0.799 3.448 0.854 ;
      RECT 3.249 0.163 3.310 0.252 ;
      RECT 3.177 0.637 3.273 0.735 ;
      RECT 2.768 0.163 3.249 0.218 ;
      RECT 3.106 0.637 3.177 0.692 ;
      RECT 3.106 0.313 3.166 0.368 ;
      RECT 3.045 0.313 3.106 0.692 ;
      RECT 3.011 0.445 3.045 0.545 ;
      RECT 2.934 0.767 2.986 0.854 ;
      RECT 2.934 0.287 2.955 0.374 ;
      RECT 2.873 0.287 2.934 0.854 ;
      RECT 2.754 0.796 2.780 0.877 ;
      RECT 2.754 0.163 2.768 0.343 ;
      RECT 2.707 0.163 2.754 0.877 ;
      RECT 2.693 0.262 2.707 0.877 ;
      RECT 2.678 0.262 2.693 0.343 ;
      RECT 2.528 0.177 2.589 0.877 ;
      RECT 2.477 0.177 2.528 0.232 ;
      RECT 2.401 0.495 2.462 0.898 ;
      RECT 1.990 0.843 2.401 0.898 ;
      RECT 2.067 0.252 2.128 0.776 ;
      RECT 1.929 0.252 1.990 0.898 ;
      RECT 1.851 0.252 1.929 0.333 ;
      RECT 1.787 0.843 1.929 0.898 ;
      RECT 1.791 0.436 1.852 0.774 ;
      RECT 1.739 0.436 1.791 0.490 ;
      RECT 1.586 0.719 1.791 0.774 ;
      RECT 1.678 0.252 1.739 0.490 ;
      RECT 1.653 0.546 1.714 0.664 ;
      RECT 1.649 0.252 1.678 0.333 ;
      RECT 1.330 0.610 1.653 0.664 ;
      RECT 1.584 0.830 1.645 1.008 ;
      RECT 0.481 0.830 1.584 0.885 ;
      RECT 1.269 0.287 1.330 0.744 ;
      RECT 1.169 0.287 1.269 0.342 ;
      RECT 0.927 0.689 1.269 0.744 ;
      RECT 0.866 0.595 0.927 0.744 ;
      RECT 0.757 0.595 0.866 0.650 ;
      RECT 0.772 0.260 0.801 0.340 ;
      RECT 0.619 0.705 0.782 0.760 ;
      RECT 0.711 0.260 0.772 0.439 ;
      RECT 0.696 0.510 0.757 0.650 ;
      RECT 0.619 0.385 0.711 0.439 ;
      RECT 0.558 0.385 0.619 0.760 ;
      RECT 0.481 0.237 0.570 0.318 ;
      RECT 0.420 0.237 0.481 0.885 ;
      RECT 0.282 0.263 0.343 0.817 ;
  END
END MXI4X2

MACRO MXI2X4
  CLASS CORE ;
  FOREIGN MXI2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.518 0.171 1.604 0.262 ;
      RECT 1.155 0.854 1.527 0.908 ;
      RECT 1.215 0.171 1.518 0.226 ;
      RECT 1.212 0.171 1.215 0.255 ;
      RECT 1.155 0.167 1.212 0.500 ;
      RECT 1.109 0.167 1.155 0.908 ;
      RECT 0.828 0.171 1.109 0.226 ;
      RECT 1.093 0.439 1.109 0.908 ;
      RECT 1.013 0.833 1.093 0.908 ;
      RECT 0.694 0.854 1.013 0.908 ;
      RECT 0.736 0.171 0.828 0.252 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.602 0.954 1.694 1.035 ;
      RECT 1.466 0.967 1.602 1.035 ;
      RECT 0.626 0.980 1.466 1.035 ;
      RECT 0.564 0.943 0.626 1.035 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.002 0.514 2.189 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.299 0.526 0.406 0.607 ;
      RECT 0.237 0.526 0.299 0.627 ;
      RECT 0.152 0.526 0.237 0.607 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.451 -0.080 2.500 0.080 ;
      RECT 2.359 -0.080 2.451 0.235 ;
      RECT 2.078 -0.080 2.359 0.080 ;
      RECT 1.986 -0.080 2.078 0.122 ;
      RECT 0.499 -0.080 1.986 0.080 ;
      RECT 0.407 -0.080 0.499 0.235 ;
      RECT 0.146 -0.080 0.407 0.080 ;
      RECT 0.054 -0.080 0.146 0.240 ;
      RECT 0.000 -0.080 0.054 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.451 1.120 2.500 1.280 ;
      RECT 2.359 0.979 2.451 1.280 ;
      RECT 2.071 1.120 2.359 1.280 ;
      RECT 1.979 0.896 2.071 1.280 ;
      RECT 0.483 1.120 1.979 1.280 ;
      RECT 0.421 0.979 0.483 1.280 ;
      RECT 0.146 1.120 0.421 1.280 ;
      RECT 0.054 0.982 0.146 1.280 ;
      RECT 0.000 1.120 0.054 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.344 0.363 2.407 0.760 ;
      RECT 2.273 0.363 2.344 0.418 ;
      RECT 2.271 0.705 2.344 0.760 ;
      RECT 2.242 0.336 2.273 0.418 ;
      RECT 2.179 0.705 2.271 0.865 ;
      RECT 2.196 0.221 2.242 0.418 ;
      RECT 2.181 0.221 2.196 0.417 ;
      RECT 2.179 0.221 2.181 0.404 ;
      RECT 1.730 0.221 2.179 0.276 ;
      RECT 1.855 0.662 1.893 0.764 ;
      RECT 1.792 0.336 1.855 0.764 ;
      RECT 1.694 0.710 1.792 0.764 ;
      RECT 1.668 0.221 1.730 0.404 ;
      RECT 1.602 0.710 1.694 0.790 ;
      RECT 1.402 0.349 1.668 0.404 ;
      RECT 1.339 0.349 1.402 0.733 ;
      RECT 1.335 0.679 1.339 0.733 ;
      RECT 1.243 0.679 1.335 0.760 ;
      RECT 0.908 0.336 1.000 0.417 ;
      RECT 0.874 0.657 0.966 0.751 ;
      RECT 0.875 0.362 0.908 0.417 ;
      RECT 0.813 0.362 0.875 0.449 ;
      RECT 0.561 0.696 0.874 0.751 ;
      RECT 0.561 0.394 0.813 0.449 ;
      RECT 0.499 0.394 0.561 0.754 ;
      RECT 0.325 0.394 0.499 0.449 ;
      RECT 0.325 0.696 0.499 0.754 ;
      RECT 0.233 0.336 0.325 0.449 ;
      RECT 0.248 0.696 0.325 0.786 ;
      RECT 0.233 0.699 0.248 0.786 ;
  END
END MXI2X4

MACRO MXI2X2
  CLASS CORE ;
  FOREIGN MXI2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.883 0.293 0.944 0.888 ;
      RECT 0.838 0.833 0.883 0.888 ;
      RECT 0.716 0.833 0.838 1.005 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.179 0.656 0.313 0.767 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.506 0.493 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.252 0.433 1.363 0.576 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.352 -0.080 1.400 0.080 ;
      RECT 1.262 -0.080 1.352 0.122 ;
      RECT 0.459 -0.080 1.262 0.080 ;
      RECT 0.369 -0.080 0.459 0.261 ;
      RECT 0.000 -0.080 0.369 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.352 1.120 1.400 1.280 ;
      RECT 1.262 0.757 1.352 1.280 ;
      RECT 0.377 1.120 1.262 1.280 ;
      RECT 0.286 0.853 0.377 1.280 ;
      RECT 0.000 1.120 0.286 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.128 0.336 1.189 0.790 ;
      RECT 1.115 0.736 1.128 0.790 ;
      RECT 1.025 0.736 1.115 0.960 ;
      RECT 1.005 0.163 1.066 0.571 ;
      RECT 0.615 0.163 1.005 0.218 ;
      RECT 0.761 0.326 0.822 0.763 ;
      RECT 0.677 0.326 0.761 0.407 ;
      RECT 0.583 0.708 0.761 0.763 ;
      RECT 0.615 0.517 0.696 0.607 ;
      RECT 0.554 0.163 0.615 0.607 ;
      RECT 0.493 0.708 0.583 1.013 ;
      RECT 0.257 0.387 0.554 0.442 ;
      RECT 0.196 0.257 0.257 0.442 ;
      RECT 0.167 0.257 0.196 0.348 ;
      RECT 0.109 0.293 0.167 0.348 ;
      RECT 0.109 0.836 0.138 0.917 ;
      RECT 0.048 0.293 0.109 0.917 ;
  END
END MXI2X2

MACRO MXI2X1
  CLASS CORE ;
  FOREIGN MXI2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.829 0.573 0.868 0.805 ;
      RECT 0.829 0.281 0.844 0.362 ;
      RECT 0.764 0.281 0.829 0.805 ;
      RECT 0.748 0.281 0.764 0.362 ;
      RECT 0.748 0.724 0.764 0.805 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.198 0.524 0.332 0.633 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.411 0.433 0.529 0.555 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.128 0.433 1.261 0.543 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.247 -0.080 1.300 0.080 ;
      RECT 1.151 -0.080 1.247 0.122 ;
      RECT 0.411 -0.080 1.151 0.080 ;
      RECT 0.315 -0.080 0.411 0.347 ;
      RECT 0.000 -0.080 0.315 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.251 1.120 1.300 1.280 ;
      RECT 1.152 1.064 1.251 1.280 ;
      RECT 0.400 1.120 1.152 1.280 ;
      RECT 0.304 0.954 0.400 1.280 ;
      RECT 0.000 1.120 0.304 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.040 0.710 1.069 0.790 ;
      RECT 1.040 0.279 1.058 0.360 ;
      RECT 0.975 0.279 1.040 0.790 ;
      RECT 0.962 0.279 0.975 0.360 ;
      RECT 0.974 0.710 0.975 0.790 ;
      RECT 0.654 0.933 0.698 1.014 ;
      RECT 0.612 0.281 0.677 0.760 ;
      RECT 0.590 0.815 0.654 1.014 ;
      RECT 0.535 0.281 0.612 0.362 ;
      RECT 0.529 0.679 0.612 0.760 ;
      RECT 0.152 0.815 0.590 0.870 ;
      RECT 0.163 0.292 0.165 0.368 ;
      RECT 0.114 0.292 0.163 0.381 ;
      RECT 0.114 0.736 0.152 0.870 ;
      RECT 0.049 0.292 0.114 0.870 ;
  END
END MXI2X1

MACRO MX4X4
  CLASS CORE ;
  FOREIGN MX4X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.887 0.320 3.988 0.900 ;
      RECT 3.865 0.320 3.887 0.424 ;
      RECT 3.865 0.657 3.887 0.900 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.430 0.579 3.513 0.660 ;
      RECT 3.369 0.579 3.430 0.894 ;
      RECT 2.938 0.839 3.369 0.894 ;
      RECT 2.837 0.839 2.938 0.919 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.024 0.951 2.085 1.033 ;
      RECT 0.757 0.951 2.024 1.006 ;
      RECT 0.643 0.951 0.757 1.014 ;
      RECT 0.630 0.951 0.643 1.027 ;
      RECT 0.618 0.960 0.630 1.027 ;
      RECT 0.528 0.960 0.618 1.040 ;
     END
  END S0

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.107 0.561 1.168 0.627 ;
      RECT 1.010 0.561 1.107 0.615 ;
      RECT 0.949 0.524 1.010 0.615 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.111 0.433 0.202 0.550 ;
      RECT 0.037 0.433 0.111 0.549 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.580 0.433 1.713 0.540 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.453 0.525 2.588 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.128 -0.080 4.200 0.080 ;
      RECT 4.038 -0.080 4.128 0.242 ;
      RECT 3.778 -0.080 4.038 0.080 ;
      RECT 3.688 -0.080 3.778 0.224 ;
      RECT 2.608 -0.080 3.688 0.080 ;
      RECT 2.518 -0.080 2.608 0.122 ;
      RECT 1.609 -0.080 2.518 0.080 ;
      RECT 1.519 -0.080 1.609 0.122 ;
      RECT 1.145 -0.080 1.519 0.080 ;
      RECT 1.055 -0.080 1.145 0.122 ;
      RECT 0.138 -0.080 1.055 0.080 ;
      RECT 0.048 -0.080 0.138 0.364 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.128 1.120 4.200 1.280 ;
      RECT 4.038 0.982 4.128 1.280 ;
      RECT 3.778 1.120 4.038 1.280 ;
      RECT 3.688 0.982 3.778 1.280 ;
      RECT 2.606 1.120 3.688 1.280 ;
      RECT 2.516 1.078 2.606 1.280 ;
      RECT 1.609 1.120 2.516 1.280 ;
      RECT 1.519 1.078 1.609 1.280 ;
      RECT 1.112 1.120 1.519 1.280 ;
      RECT 1.022 1.078 1.112 1.280 ;
      RECT 0.138 1.120 1.022 1.280 ;
      RECT 0.048 0.757 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.682 0.299 3.743 0.787 ;
      RECT 3.538 0.299 3.682 0.354 ;
      RECT 3.554 0.732 3.682 0.787 ;
      RECT 3.529 0.408 3.615 0.508 ;
      RECT 3.493 0.732 3.554 1.042 ;
      RECT 3.448 0.157 3.538 0.354 ;
      RECT 3.317 0.437 3.529 0.492 ;
      RECT 2.744 0.987 3.493 1.042 ;
      RECT 3.239 0.194 3.317 0.492 ;
      RECT 3.227 0.194 3.239 0.762 ;
      RECT 3.178 0.437 3.227 0.762 ;
      RECT 3.134 0.681 3.178 0.762 ;
      RECT 3.077 0.200 3.106 0.402 ;
      RECT 3.019 0.200 3.077 0.592 ;
      RECT 3.019 0.681 3.033 0.762 ;
      RECT 3.016 0.200 3.019 0.762 ;
      RECT 2.203 0.200 3.016 0.255 ;
      RECT 2.958 0.537 3.016 0.762 ;
      RECT 2.943 0.681 2.958 0.762 ;
      RECT 2.795 0.336 2.950 0.417 ;
      RECT 2.795 0.688 2.809 0.769 ;
      RECT 2.734 0.336 2.795 0.769 ;
      RECT 2.683 0.939 2.744 1.042 ;
      RECT 2.719 0.336 2.734 0.417 ;
      RECT 2.719 0.688 2.734 0.769 ;
      RECT 2.231 0.939 2.683 0.994 ;
      RECT 2.370 0.317 2.400 0.398 ;
      RECT 2.370 0.692 2.400 0.885 ;
      RECT 2.309 0.317 2.370 0.885 ;
      RECT 2.170 0.842 2.231 0.994 ;
      RECT 2.154 0.200 2.203 0.310 ;
      RECT 1.567 0.842 2.170 0.896 ;
      RECT 2.154 0.679 2.169 0.760 ;
      RECT 2.101 0.200 2.154 0.760 ;
      RECT 2.093 0.206 2.101 0.760 ;
      RECT 2.079 0.679 2.093 0.760 ;
      RECT 1.955 0.329 2.016 0.773 ;
      RECT 1.819 0.329 1.955 0.410 ;
      RECT 1.811 0.718 1.955 0.773 ;
      RECT 1.823 0.150 1.909 0.205 ;
      RECT 1.879 0.526 1.893 0.607 ;
      RECT 1.803 0.526 1.879 0.650 ;
      RECT 1.762 0.150 1.823 0.261 ;
      RECT 1.721 0.705 1.811 0.786 ;
      RECT 1.348 0.595 1.803 0.650 ;
      RECT 0.846 0.206 1.762 0.261 ;
      RECT 1.506 0.825 1.567 0.896 ;
      RECT 1.175 0.825 1.506 0.880 ;
      RECT 1.328 0.346 1.348 0.650 ;
      RECT 1.267 0.346 1.328 0.770 ;
      RECT 1.252 0.346 1.267 0.411 ;
      RECT 1.238 0.689 1.267 0.770 ;
      RECT 0.871 0.346 1.252 0.401 ;
      RECT 1.114 0.814 1.175 0.880 ;
      RECT 0.520 0.814 1.114 0.869 ;
      RECT 0.817 0.679 0.907 0.760 ;
      RECT 0.810 0.346 0.871 0.605 ;
      RECT 0.756 0.171 0.846 0.261 ;
      RECT 0.671 0.692 0.817 0.746 ;
      RECT 0.734 0.524 0.810 0.605 ;
      RECT 0.671 0.325 0.748 0.406 ;
      RECT 0.610 0.325 0.671 0.746 ;
      RECT 0.510 0.186 0.521 0.379 ;
      RECT 0.510 0.814 0.520 0.895 ;
      RECT 0.449 0.186 0.510 0.895 ;
      RECT 0.431 0.186 0.449 0.379 ;
      RECT 0.430 0.814 0.449 0.895 ;
      RECT 0.268 0.186 0.329 0.965 ;
      RECT 0.239 0.186 0.268 0.379 ;
      RECT 0.239 0.742 0.268 0.965 ;
  END
END MX4X4

MACRO MX4X2
  CLASS CORE ;
  FOREIGN MX4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.906 0.706 3.943 0.761 ;
      RECT 3.846 0.180 3.906 1.006 ;
      RECT 3.817 0.180 3.846 0.373 ;
      RECT 3.817 0.701 3.846 1.006 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.408 0.579 3.491 0.660 ;
      RECT 3.348 0.579 3.408 0.894 ;
      RECT 2.920 0.839 3.348 0.894 ;
      RECT 2.819 0.839 2.920 0.919 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.012 0.951 2.072 1.033 ;
      RECT 0.752 0.951 2.012 1.006 ;
      RECT 0.639 0.951 0.752 1.014 ;
      RECT 0.626 0.951 0.639 1.027 ;
      RECT 0.614 0.960 0.626 1.027 ;
      RECT 0.524 0.960 0.614 1.040 ;
     END
  END S0

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.100 0.561 1.161 0.627 ;
      RECT 1.004 0.561 1.100 0.615 ;
      RECT 0.943 0.524 1.004 0.615 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.111 0.433 0.200 0.550 ;
      RECT 0.037 0.433 0.111 0.549 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.570 0.433 1.702 0.540 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.437 0.525 2.572 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.701 -0.080 4.000 0.080 ;
      RECT 3.611 -0.080 3.701 0.210 ;
      RECT 2.592 -0.080 3.611 0.080 ;
      RECT 2.502 -0.080 2.592 0.122 ;
      RECT 1.599 -0.080 2.502 0.080 ;
      RECT 1.510 -0.080 1.599 0.122 ;
      RECT 1.138 -0.080 1.510 0.080 ;
      RECT 1.049 -0.080 1.138 0.122 ;
      RECT 0.137 -0.080 1.049 0.080 ;
      RECT 0.047 -0.080 0.137 0.364 ;
      RECT 0.000 -0.080 0.047 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.701 1.120 4.000 1.280 ;
      RECT 3.611 0.877 3.701 1.280 ;
      RECT 2.590 1.120 3.611 1.280 ;
      RECT 2.501 1.078 2.590 1.280 ;
      RECT 1.599 1.120 2.501 1.280 ;
      RECT 1.510 1.078 1.599 1.280 ;
      RECT 1.105 1.120 1.510 1.280 ;
      RECT 1.016 1.078 1.105 1.280 ;
      RECT 0.137 1.120 1.016 1.280 ;
      RECT 0.047 0.757 0.137 1.280 ;
      RECT 0.000 1.120 0.047 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.659 0.295 3.719 0.787 ;
      RECT 3.516 0.295 3.659 0.350 ;
      RECT 3.532 0.732 3.659 0.787 ;
      RECT 3.507 0.408 3.593 0.508 ;
      RECT 3.472 0.732 3.532 1.042 ;
      RECT 3.427 0.157 3.516 0.350 ;
      RECT 3.296 0.437 3.507 0.492 ;
      RECT 2.727 0.987 3.472 1.042 ;
      RECT 3.207 0.194 3.296 0.492 ;
      RECT 3.204 0.437 3.207 0.492 ;
      RECT 3.144 0.437 3.204 0.762 ;
      RECT 3.115 0.681 3.144 0.762 ;
      RECT 3.058 0.200 3.087 0.402 ;
      RECT 3.000 0.200 3.058 0.592 ;
      RECT 3.000 0.681 3.014 0.762 ;
      RECT 2.997 0.200 3.000 0.762 ;
      RECT 2.190 0.200 2.997 0.255 ;
      RECT 2.939 0.537 2.997 0.762 ;
      RECT 2.925 0.681 2.939 0.762 ;
      RECT 2.777 0.336 2.931 0.417 ;
      RECT 2.777 0.688 2.792 0.769 ;
      RECT 2.717 0.336 2.777 0.769 ;
      RECT 2.667 0.939 2.727 1.042 ;
      RECT 2.702 0.336 2.717 0.417 ;
      RECT 2.702 0.688 2.717 0.769 ;
      RECT 2.217 0.939 2.667 0.994 ;
      RECT 2.356 0.317 2.385 0.398 ;
      RECT 2.356 0.692 2.385 0.885 ;
      RECT 2.295 0.317 2.356 0.885 ;
      RECT 2.157 0.842 2.217 0.994 ;
      RECT 2.141 0.200 2.190 0.310 ;
      RECT 1.557 0.842 2.157 0.896 ;
      RECT 2.141 0.679 2.155 0.760 ;
      RECT 2.088 0.200 2.141 0.760 ;
      RECT 2.080 0.206 2.088 0.760 ;
      RECT 2.066 0.679 2.080 0.760 ;
      RECT 1.943 0.329 2.004 0.773 ;
      RECT 1.808 0.329 1.943 0.410 ;
      RECT 1.800 0.718 1.943 0.773 ;
      RECT 1.812 0.150 1.897 0.205 ;
      RECT 1.867 0.526 1.881 0.607 ;
      RECT 1.792 0.526 1.867 0.650 ;
      RECT 1.751 0.150 1.812 0.261 ;
      RECT 1.710 0.705 1.800 0.786 ;
      RECT 1.340 0.595 1.792 0.650 ;
      RECT 0.841 0.206 1.751 0.261 ;
      RECT 1.497 0.825 1.557 0.896 ;
      RECT 1.167 0.825 1.497 0.880 ;
      RECT 1.320 0.346 1.340 0.650 ;
      RECT 1.260 0.346 1.320 0.770 ;
      RECT 1.244 0.346 1.260 0.411 ;
      RECT 1.231 0.689 1.260 0.770 ;
      RECT 0.866 0.346 1.244 0.401 ;
      RECT 1.107 0.814 1.167 0.880 ;
      RECT 0.516 0.814 1.107 0.869 ;
      RECT 0.812 0.679 0.901 0.760 ;
      RECT 0.805 0.346 0.866 0.605 ;
      RECT 0.751 0.171 0.841 0.261 ;
      RECT 0.667 0.692 0.812 0.746 ;
      RECT 0.730 0.524 0.805 0.605 ;
      RECT 0.667 0.325 0.743 0.406 ;
      RECT 0.606 0.325 0.667 0.746 ;
      RECT 0.507 0.186 0.518 0.379 ;
      RECT 0.507 0.814 0.516 0.895 ;
      RECT 0.447 0.186 0.507 0.895 ;
      RECT 0.428 0.186 0.447 0.379 ;
      RECT 0.427 0.814 0.447 0.895 ;
      RECT 0.266 0.186 0.327 0.965 ;
      RECT 0.237 0.186 0.266 0.379 ;
      RECT 0.237 0.742 0.266 0.965 ;
  END
END MX4X2

MACRO MX2X4
  CLASS CORE ;
  FOREIGN MX2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.478 0.167 1.582 0.798 ;
      RECT 1.424 0.707 1.478 0.798 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.266 0.700 0.502 0.767 ;
      RECT 0.170 0.677 0.266 0.767 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.235 0.421 0.413 0.512 ;
      RECT 0.218 0.433 0.235 0.512 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.118 0.433 1.261 0.533 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.748 -0.080 1.800 0.080 ;
      RECT 1.655 -0.080 1.748 0.211 ;
      RECT 1.372 -0.080 1.655 0.080 ;
      RECT 1.279 -0.080 1.372 0.211 ;
      RECT 0.398 -0.080 1.279 0.080 ;
      RECT 0.305 -0.080 0.398 0.352 ;
      RECT 0.000 -0.080 0.305 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.745 1.120 1.800 1.280 ;
      RECT 1.653 1.078 1.745 1.280 ;
      RECT 1.320 1.120 1.653 1.280 ;
      RECT 1.227 0.986 1.320 1.280 ;
      RECT 0.355 1.120 1.227 1.280 ;
      RECT 0.262 0.855 0.355 1.280 ;
      RECT 0.000 1.120 0.262 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.729 0.495 1.744 0.576 ;
      RECT 1.666 0.495 1.729 0.914 ;
      RECT 1.651 0.495 1.666 0.576 ;
      RECT 0.919 0.860 1.666 0.914 ;
      RECT 1.324 0.313 1.387 0.651 ;
      RECT 1.107 0.313 1.324 0.368 ;
      RECT 1.094 0.596 1.324 0.651 ;
      RECT 1.031 0.596 1.094 0.788 ;
      RECT 0.982 0.161 1.045 0.507 ;
      RECT 1.001 0.707 1.031 0.788 ;
      RECT 0.556 0.161 0.982 0.215 ;
      RECT 0.856 0.290 0.919 0.914 ;
      RECT 0.712 0.833 0.856 0.914 ;
      RECT 0.709 0.290 0.772 0.758 ;
      RECT 0.620 0.290 0.709 0.371 ;
      RECT 0.648 0.704 0.709 0.758 ;
      RECT 0.585 0.704 0.648 0.892 ;
      RECT 0.556 0.475 0.642 0.557 ;
      RECT 0.567 0.837 0.585 0.892 ;
      RECT 0.475 0.837 0.567 0.918 ;
      RECT 0.494 0.161 0.556 0.621 ;
      RECT 0.108 0.567 0.494 0.621 ;
      RECT 0.108 0.293 0.147 0.374 ;
      RECT 0.108 0.840 0.147 0.921 ;
      RECT 0.045 0.293 0.108 0.921 ;
  END
END MX2X4

MACRO MX2X2
  CLASS CORE ;
  FOREIGN MX2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.494 0.194 1.556 0.977 ;
      RECT 1.480 0.194 1.494 0.439 ;
      RECT 1.446 0.700 1.494 0.977 ;
      RECT 1.461 0.194 1.480 0.395 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.302 0.706 0.475 0.761 ;
      RECT 0.225 0.706 0.302 0.795 ;
      RECT 0.210 0.714 0.225 0.795 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.215 0.526 0.387 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.285 0.306 1.364 0.361 ;
      RECT 1.222 0.306 1.285 0.367 ;
      RECT 1.160 0.306 1.222 0.575 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 -0.080 1.600 0.080 ;
      RECT 1.244 -0.080 1.336 0.223 ;
      RECT 0.407 -0.080 1.244 0.080 ;
      RECT 0.315 -0.080 0.407 0.296 ;
      RECT 0.000 -0.080 0.315 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.323 1.120 1.600 1.280 ;
      RECT 1.231 1.078 1.323 1.280 ;
      RECT 0.407 1.120 1.231 1.280 ;
      RECT 0.315 0.890 0.407 1.280 ;
      RECT 0.000 1.120 0.315 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.385 0.485 1.415 0.595 ;
      RECT 1.323 0.485 1.385 0.994 ;
      RECT 0.941 0.939 1.323 0.994 ;
      RECT 1.020 0.279 1.081 0.858 ;
      RECT 0.879 0.267 0.941 0.994 ;
      RECT 0.843 0.267 0.879 0.321 ;
      RECT 0.770 0.836 0.879 0.917 ;
      RECT 0.752 0.240 0.843 0.321 ;
      RECT 0.739 0.396 0.801 0.761 ;
      RECT 0.667 0.396 0.739 0.451 ;
      RECT 0.642 0.706 0.739 0.761 ;
      RECT 0.605 0.190 0.667 0.451 ;
      RECT 0.599 0.520 0.661 0.606 ;
      RECT 0.580 0.706 0.642 0.915 ;
      RECT 0.547 0.190 0.605 0.245 ;
      RECT 0.527 0.520 0.599 0.575 ;
      RECT 0.465 0.370 0.527 0.575 ;
      RECT 0.140 0.370 0.465 0.425 ;
      RECT 0.125 0.858 0.145 0.939 ;
      RECT 0.125 0.348 0.140 0.429 ;
      RECT 0.063 0.348 0.125 0.939 ;
      RECT 0.048 0.348 0.063 0.429 ;
      RECT 0.054 0.858 0.063 0.939 ;
  END
END MX2X2

MACRO MX2X1
  CLASS CORE ;
  FOREIGN MX2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.302 0.268 1.363 0.946 ;
      RECT 1.250 0.268 1.302 0.379 ;
      RECT 1.198 0.754 1.302 0.946 ;
      RECT 1.248 0.268 1.250 0.361 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.944 0.188 1.033 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.688 0.488 0.767 ;
      RECT 0.292 0.635 0.387 0.767 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.000 0.433 1.188 0.527 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.139 -0.080 1.400 0.080 ;
      RECT 1.049 -0.080 1.139 0.122 ;
      RECT 0.349 -0.080 1.049 0.080 ;
      RECT 0.349 0.291 0.351 0.342 ;
      RECT 0.264 -0.080 0.349 0.342 ;
      RECT 0.000 -0.080 0.264 0.080 ;
      RECT 0.261 0.291 0.264 0.342 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.140 1.120 1.400 1.280 ;
      RECT 1.050 1.078 1.140 1.280 ;
      RECT 0.339 1.120 1.050 1.280 ;
      RECT 0.249 0.852 0.339 1.280 ;
      RECT 0.000 1.120 0.249 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.103 0.615 1.193 0.696 ;
      RECT 1.096 0.621 1.103 0.696 ;
      RECT 1.035 0.621 1.096 0.968 ;
      RECT 0.793 0.913 1.035 0.968 ;
      RECT 0.862 0.269 0.923 0.838 ;
      RECT 0.732 0.280 0.793 0.968 ;
      RECT 0.654 0.280 0.732 0.335 ;
      RECT 0.671 0.789 0.732 0.882 ;
      RECT 0.610 0.393 0.671 0.720 ;
      RECT 0.553 0.393 0.610 0.448 ;
      RECT 0.549 0.665 0.610 0.887 ;
      RECT 0.492 0.269 0.553 0.448 ;
      RECT 0.440 0.832 0.549 0.887 ;
      RECT 0.460 0.508 0.546 0.599 ;
      RECT 0.463 0.269 0.492 0.350 ;
      RECT 0.123 0.524 0.460 0.579 ;
      RECT 0.123 0.276 0.138 0.357 ;
      RECT 0.123 0.752 0.138 0.833 ;
      RECT 0.062 0.276 0.123 0.833 ;
      RECT 0.048 0.276 0.062 0.357 ;
      RECT 0.048 0.752 0.062 0.833 ;
  END
END MX2X1

MACRO INVXL
  CLASS CORE ;
  FOREIGN INVXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.312 0.567 0.358 0.768 ;
      RECT 0.312 0.321 0.339 0.439 ;
      RECT 0.242 0.321 0.312 0.768 ;
      RECT 0.236 0.321 0.242 0.439 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.158 0.598 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.300 -0.080 0.400 0.080 ;
      RECT 0.055 -0.080 0.300 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.258 1.120 0.400 1.280 ;
      RECT 0.258 0.925 0.329 0.975 ;
      RECT 0.155 0.925 0.258 1.280 ;
      RECT 0.083 0.925 0.155 0.975 ;
      RECT 0.000 1.120 0.155 1.280 ;
     END
  END VDD
END INVXL

MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.878 0.419 1.040 0.767 ;
      RECT 0.857 0.361 0.878 0.767 ;
      RECT 0.811 0.361 0.857 0.780 ;
      RECT 0.610 0.307 0.811 0.812 ;
      RECT 0.589 0.307 0.610 0.433 ;
      RECT 0.217 0.698 0.610 0.812 ;
      RECT 0.217 0.307 0.589 0.421 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.150 0.487 0.376 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.043 -0.080 1.100 0.080 ;
      RECT 0.818 -0.080 1.043 0.122 ;
      RECT 0.533 -0.080 0.818 0.080 ;
      RECT 0.439 -0.080 0.533 0.214 ;
      RECT 0.156 -0.080 0.439 0.080 ;
      RECT 0.061 -0.080 0.156 0.122 ;
      RECT 0.000 -0.080 0.061 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 1.120 1.100 1.280 ;
      RECT 0.922 1.078 1.050 1.280 ;
      RECT 0.828 0.917 0.922 1.280 ;
      RECT 0.532 1.120 0.828 1.280 ;
      RECT 0.438 0.917 0.532 1.280 ;
      RECT 0.144 1.120 0.438 1.280 ;
      RECT 0.050 0.917 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
END INVX8

MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.251 0.194 0.341 1.010 ;
      RECT 0.212 0.433 0.251 0.767 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.446 0.138 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.542 -0.080 0.700 0.080 ;
      RECT 0.452 -0.080 0.542 0.372 ;
      RECT 0.138 -0.080 0.452 0.080 ;
      RECT 0.048 -0.080 0.138 0.372 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.542 1.120 0.700 1.280 ;
      RECT 0.452 0.720 0.542 1.280 ;
      RECT 0.138 1.120 0.452 1.280 ;
      RECT 0.048 0.720 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
END INVX4

MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.183 0.558 0.715 ;
      RECT 0.442 0.183 0.488 0.376 ;
      RECT 0.465 0.627 0.488 0.715 ;
      RECT 0.327 0.661 0.465 0.715 ;
      RECT 0.224 0.661 0.327 0.854 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.150 0.433 0.395 0.574 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.267 -0.080 0.600 0.080 ;
      RECT 0.164 -0.080 0.267 0.361 ;
      RECT 0.000 -0.080 0.164 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.497 1.120 0.600 1.280 ;
      RECT 0.495 1.078 0.497 1.280 ;
      RECT 0.395 1.064 0.495 1.280 ;
      RECT 0.394 1.078 0.395 1.280 ;
      RECT 0.000 1.120 0.394 1.280 ;
     END
  END VDD
END INVX2

MACRO INVX20
  CLASS CORE ;
  FOREIGN INVX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.836 0.285 3.243 0.914 ;
      RECT 2.733 0.285 2.836 0.448 ;
      RECT 2.693 0.712 2.836 0.874 ;
      RECT 1.899 0.286 2.733 0.448 ;
      RECT 2.549 0.696 2.693 0.889 ;
      RECT 2.320 0.712 2.549 0.874 ;
      RECT 2.201 0.696 2.320 0.889 ;
      RECT 1.967 0.712 2.201 0.874 ;
      RECT 1.854 0.696 1.967 0.889 ;
      RECT 1.809 0.285 1.899 0.448 ;
      RECT 1.620 0.712 1.854 0.874 ;
      RECT 1.480 0.285 1.809 0.446 ;
      RECT 1.480 0.696 1.620 0.889 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.211 0.500 0.330 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.246 -0.080 3.300 0.080 ;
      RECT 3.157 -0.080 3.246 0.122 ;
      RECT 2.882 -0.080 3.157 0.080 ;
      RECT 2.792 -0.080 2.882 0.122 ;
      RECT 2.508 -0.080 2.792 0.080 ;
      RECT 2.418 -0.080 2.508 0.122 ;
      RECT 2.132 -0.080 2.418 0.080 ;
      RECT 2.042 -0.080 2.132 0.122 ;
      RECT 1.758 -0.080 2.042 0.080 ;
      RECT 1.668 -0.080 1.758 0.122 ;
      RECT 1.391 -0.080 1.668 0.080 ;
      RECT 1.301 -0.080 1.391 0.122 ;
      RECT 1.011 -0.080 1.301 0.080 ;
      RECT 0.921 -0.080 1.011 0.228 ;
      RECT 0.636 -0.080 0.921 0.080 ;
      RECT 0.546 -0.080 0.636 0.228 ;
      RECT 0.264 -0.080 0.546 0.080 ;
      RECT 0.175 -0.080 0.264 0.386 ;
      RECT 0.000 -0.080 0.175 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.246 1.120 3.300 1.280 ;
      RECT 3.157 1.078 3.246 1.280 ;
      RECT 2.882 1.120 3.157 1.280 ;
      RECT 2.792 1.078 2.882 1.280 ;
      RECT 2.508 1.120 2.792 1.280 ;
      RECT 2.418 1.078 2.508 1.280 ;
      RECT 2.130 1.120 2.418 1.280 ;
      RECT 2.041 1.078 2.130 1.280 ;
      RECT 1.757 1.120 2.041 1.280 ;
      RECT 1.667 1.078 1.757 1.280 ;
      RECT 1.384 1.120 1.667 1.280 ;
      RECT 1.295 1.078 1.384 1.280 ;
      RECT 1.009 1.120 1.295 1.280 ;
      RECT 0.920 0.982 1.009 1.280 ;
      RECT 0.622 1.120 0.920 1.280 ;
      RECT 0.533 0.989 0.622 1.280 ;
      RECT 0.264 1.120 0.533 1.280 ;
      RECT 0.175 0.741 0.264 1.280 ;
      RECT 0.000 1.120 0.175 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.425 0.521 2.751 0.602 ;
      RECT 1.268 0.526 1.425 0.598 ;
      RECT 1.189 0.338 1.268 0.889 ;
      RECT 0.734 0.338 1.189 0.419 ;
      RECT 0.733 0.696 1.189 0.889 ;
      RECT 0.653 0.500 1.113 0.581 ;
      RECT 0.467 0.513 0.653 0.568 ;
      RECT 0.407 0.338 0.467 0.789 ;
      RECT 0.378 0.338 0.407 0.419 ;
      RECT 0.378 0.708 0.407 0.789 ;
  END
END INVX20

MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.323 0.564 0.358 0.848 ;
      RECT 0.253 0.321 0.323 0.848 ;
      RECT 0.242 0.564 0.253 0.848 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.173 0.568 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 -0.080 0.400 0.080 ;
      RECT 0.055 -0.080 0.158 0.122 ;
      RECT 0.000 -0.080 0.055 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 1.120 0.400 1.280 ;
      RECT 0.055 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.055 1.280 ;
     END
  END VDD
END INVX1

MACRO INVX16
  CLASS CORE ;
  FOREIGN INVX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.528 0.286 2.943 0.914 ;
      RECT 1.929 0.286 2.528 0.448 ;
      RECT 2.357 0.712 2.528 0.874 ;
      RECT 2.237 0.696 2.357 0.889 ;
      RECT 1.999 0.712 2.237 0.874 ;
      RECT 1.884 0.696 1.999 0.889 ;
      RECT 1.838 0.285 1.929 0.448 ;
      RECT 1.646 0.712 1.884 0.874 ;
      RECT 1.504 0.285 1.838 0.446 ;
      RECT 1.504 0.696 1.646 0.889 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.214 0.500 0.336 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.928 -0.080 3.000 0.080 ;
      RECT 2.837 -0.080 2.928 0.122 ;
      RECT 2.548 -0.080 2.837 0.080 ;
      RECT 2.457 -0.080 2.548 0.122 ;
      RECT 2.166 -0.080 2.457 0.080 ;
      RECT 2.075 -0.080 2.166 0.122 ;
      RECT 1.785 -0.080 2.075 0.080 ;
      RECT 1.694 -0.080 1.785 0.122 ;
      RECT 1.413 -0.080 1.694 0.080 ;
      RECT 1.322 -0.080 1.413 0.122 ;
      RECT 1.027 -0.080 1.322 0.080 ;
      RECT 0.936 -0.080 1.027 0.228 ;
      RECT 0.646 -0.080 0.936 0.080 ;
      RECT 0.555 -0.080 0.646 0.228 ;
      RECT 0.258 -0.080 0.555 0.080 ;
      RECT 0.167 -0.080 0.258 0.409 ;
      RECT 0.000 -0.080 0.167 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.928 1.120 3.000 1.280 ;
      RECT 2.837 1.078 2.928 1.280 ;
      RECT 2.548 1.120 2.837 1.280 ;
      RECT 2.457 1.078 2.548 1.280 ;
      RECT 2.164 1.120 2.457 1.280 ;
      RECT 2.074 1.078 2.164 1.280 ;
      RECT 1.785 1.120 2.074 1.280 ;
      RECT 1.694 1.078 1.785 1.280 ;
      RECT 1.409 1.120 1.694 1.280 ;
      RECT 1.318 1.078 1.409 1.280 ;
      RECT 1.025 1.120 1.318 1.280 ;
      RECT 0.934 0.982 1.025 1.280 ;
      RECT 0.632 1.120 0.934 1.280 ;
      RECT 0.541 0.989 0.632 1.280 ;
      RECT 0.258 1.120 0.541 1.280 ;
      RECT 0.167 0.741 0.258 1.280 ;
      RECT 0.000 1.120 0.167 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.476 0.521 2.447 0.602 ;
      RECT 1.289 0.526 1.476 0.598 ;
      RECT 1.209 0.338 1.289 0.768 ;
      RECT 0.746 0.338 1.209 0.419 ;
      RECT 1.199 0.696 1.209 0.768 ;
      RECT 1.108 0.696 1.199 0.889 ;
      RECT 0.663 0.500 1.131 0.581 ;
      RECT 0.836 0.696 1.108 0.777 ;
      RECT 0.745 0.696 0.836 0.889 ;
      RECT 0.475 0.513 0.663 0.568 ;
      RECT 0.413 0.338 0.475 0.789 ;
      RECT 0.384 0.338 0.413 0.419 ;
      RECT 0.384 0.708 0.413 0.789 ;
  END
END INVX16

MACRO INVX12
  CLASS CORE ;
  FOREIGN INVX12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.827 0.286 2.242 0.914 ;
      RECT 1.155 0.286 1.827 0.448 ;
      RECT 1.807 0.626 1.827 0.914 ;
      RECT 1.154 0.676 1.807 0.914 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.139 0.507 0.231 0.588 ;
      RECT 0.119 0.533 0.139 0.588 ;
      RECT 0.058 0.533 0.119 0.627 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.249 -0.080 2.300 0.080 ;
      RECT 2.158 -0.080 2.249 0.199 ;
      RECT 1.868 -0.080 2.158 0.080 ;
      RECT 1.777 -0.080 1.868 0.199 ;
      RECT 1.484 -0.080 1.777 0.080 ;
      RECT 1.393 -0.080 1.484 0.199 ;
      RECT 0.745 -0.080 1.393 0.080 ;
      RECT 0.654 -0.080 0.745 0.122 ;
      RECT 0.374 -0.080 0.654 0.080 ;
      RECT 0.283 -0.080 0.374 0.237 ;
      RECT 0.000 -0.080 0.283 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.252 1.120 2.300 1.280 ;
      RECT 2.161 0.989 2.252 1.280 ;
      RECT 1.868 1.120 2.161 1.280 ;
      RECT 1.777 0.989 1.868 1.280 ;
      RECT 1.484 1.120 1.777 1.280 ;
      RECT 1.393 0.989 1.484 1.280 ;
      RECT 1.110 1.120 1.393 1.280 ;
      RECT 1.017 1.065 1.110 1.280 ;
      RECT 0.359 1.120 1.017 1.280 ;
      RECT 0.268 1.078 0.359 1.280 ;
      RECT 0.000 1.120 0.268 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.936 0.521 1.745 0.602 ;
      RECT 0.855 0.338 0.936 0.767 ;
      RECT 0.470 0.338 0.855 0.419 ;
      RECT 0.562 0.686 0.855 0.767 ;
      RECT 0.379 0.500 0.713 0.581 ;
      RECT 0.470 0.686 0.562 0.888 ;
      RECT 0.318 0.343 0.379 0.770 ;
      RECT 0.145 0.343 0.318 0.398 ;
      RECT 0.139 0.715 0.318 0.770 ;
      RECT 0.054 0.343 0.145 0.424 ;
      RECT 0.048 0.689 0.139 0.770 ;
  END
END INVX12

MACRO DFFRHQX1
  CLASS CORE ;
  FOREIGN DFFRHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.099 0.693 3.310 0.776 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.639 0.296 3.643 0.761 ;
      RECT 3.581 0.296 3.639 1.021 ;
      RECT 3.356 0.296 3.581 0.351 ;
      RECT 3.561 0.706 3.581 1.021 ;
      RECT 3.548 0.829 3.561 1.021 ;
      RECT 3.294 0.174 3.356 0.351 ;
      RECT 3.265 0.174 3.294 0.255 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.431 0.306 0.471 0.361 ;
      RECT 0.431 0.431 0.432 0.512 ;
      RECT 0.370 0.306 0.431 0.512 ;
      RECT 0.342 0.431 0.370 0.512 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.240 0.573 0.295 0.633 ;
      RECT 0.155 0.517 0.240 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.548 -0.080 3.700 0.080 ;
      RECT 3.457 -0.080 3.548 0.211 ;
      RECT 3.151 -0.080 3.457 0.080 ;
      RECT 2.900 -0.080 3.151 0.122 ;
      RECT 2.596 -0.080 2.900 0.080 ;
      RECT 2.505 -0.080 2.596 0.122 ;
      RECT 1.814 -0.080 2.505 0.080 ;
      RECT 1.723 -0.080 1.814 0.254 ;
      RECT 1.073 -0.080 1.723 0.080 ;
      RECT 0.982 -0.080 1.073 0.327 ;
      RECT 0.346 -0.080 0.982 0.080 ;
      RECT 0.255 -0.080 0.346 0.234 ;
      RECT 0.000 -0.080 0.255 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.297 1.120 3.700 1.280 ;
      RECT 3.206 0.853 3.297 1.280 ;
      RECT 2.694 1.120 3.206 1.280 ;
      RECT 2.583 1.078 2.694 1.280 ;
      RECT 1.926 1.120 2.583 1.280 ;
      RECT 1.815 1.078 1.926 1.280 ;
      RECT 1.078 1.120 1.815 1.280 ;
      RECT 0.988 0.963 1.078 1.280 ;
      RECT 0.422 1.120 0.988 1.280 ;
      RECT 0.331 0.920 0.422 1.280 ;
      RECT 0.000 1.120 0.331 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.420 0.407 3.510 0.488 ;
      RECT 3.139 0.407 3.420 0.462 ;
      RECT 3.001 0.583 3.388 0.638 ;
      RECT 3.078 0.206 3.139 0.462 ;
      RECT 3.013 0.952 3.103 1.033 ;
      RECT 2.692 0.206 3.078 0.261 ;
      RECT 2.858 0.952 3.013 1.007 ;
      RECT 2.916 0.327 3.001 0.638 ;
      RECT 2.900 0.327 2.916 0.408 ;
      RECT 2.858 0.526 2.916 0.638 ;
      RECT 2.826 0.526 2.858 1.007 ;
      RECT 2.796 0.573 2.826 1.007 ;
      RECT 2.795 0.939 2.796 1.007 ;
      RECT 1.544 0.939 2.795 0.994 ;
      RECT 2.686 0.336 2.776 0.417 ;
      RECT 2.593 0.206 2.692 0.273 ;
      RECT 2.680 0.362 2.686 0.417 ;
      RECT 2.619 0.362 2.680 0.833 ;
      RECT 2.568 0.614 2.619 0.833 ;
      RECT 2.463 0.206 2.593 0.261 ;
      RECT 2.524 0.614 2.568 0.698 ;
      RECT 2.401 0.206 2.463 0.857 ;
      RECT 2.217 0.206 2.401 0.263 ;
      RECT 2.315 0.802 2.401 0.857 ;
      RECT 2.264 0.382 2.316 0.463 ;
      RECT 2.224 0.802 2.315 0.883 ;
      RECT 2.225 0.382 2.264 0.727 ;
      RECT 2.202 0.383 2.225 0.727 ;
      RECT 2.156 0.206 2.217 0.304 ;
      RECT 2.122 0.380 2.141 0.882 ;
      RECT 2.086 0.380 2.122 0.883 ;
      RECT 2.080 0.267 2.086 0.883 ;
      RECT 2.025 0.267 2.080 0.435 ;
      RECT 2.032 0.802 2.080 0.883 ;
      RECT 2.018 0.267 2.025 0.321 ;
      RECT 1.927 0.240 2.018 0.321 ;
      RECT 1.958 0.548 2.018 0.644 ;
      RECT 1.897 0.390 1.958 0.852 ;
      RECT 1.682 0.390 1.897 0.445 ;
      RECT 1.770 0.798 1.897 0.852 ;
      RECT 1.771 0.518 1.833 0.694 ;
      RECT 1.299 0.518 1.771 0.573 ;
      RECT 1.679 0.798 1.770 0.879 ;
      RECT 1.646 0.364 1.682 0.445 ;
      RECT 1.584 0.176 1.646 0.445 ;
      RECT 1.244 0.176 1.584 0.231 ;
      RECT 1.483 0.627 1.544 0.994 ;
      RECT 1.420 0.627 1.483 0.708 ;
      RECT 1.247 0.424 1.299 0.876 ;
      RECT 1.237 0.398 1.247 0.876 ;
      RECT 1.153 0.150 1.244 0.231 ;
      RECT 1.156 0.398 1.237 0.479 ;
      RECT 1.177 0.795 1.237 0.876 ;
      RECT 1.085 0.614 1.176 0.701 ;
      RECT 0.969 0.424 1.156 0.479 ;
      RECT 0.773 0.646 1.085 0.701 ;
      RECT 0.908 0.424 0.969 0.564 ;
      RECT 0.878 0.483 0.908 0.564 ;
      RECT 0.755 0.890 0.846 0.971 ;
      RECT 0.761 0.249 0.773 0.701 ;
      RECT 0.711 0.249 0.761 0.792 ;
      RECT 0.609 0.890 0.755 0.945 ;
      RECT 0.710 0.249 0.711 0.304 ;
      RECT 0.698 0.646 0.711 0.792 ;
      RECT 0.619 0.223 0.710 0.304 ;
      RECT 0.670 0.711 0.698 0.792 ;
      RECT 0.609 0.436 0.623 0.517 ;
      RECT 0.547 0.436 0.609 0.945 ;
      RECT 0.533 0.436 0.547 0.517 ;
      RECT 0.208 0.688 0.547 0.743 ;
      RECT 0.117 0.688 0.208 0.769 ;
      RECT 0.093 0.305 0.139 0.386 ;
      RECT 0.093 0.688 0.117 0.743 ;
      RECT 0.032 0.305 0.093 0.743 ;
  END
END DFFRHQX1

MACRO CLKINVX8
  CLASS CORE ;
  FOREIGN CLKINVX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.878 0.433 1.040 0.767 ;
      RECT 0.857 0.360 0.878 0.767 ;
      RECT 0.800 0.360 0.857 0.780 ;
      RECT 0.610 0.294 0.800 0.812 ;
      RECT 0.589 0.294 0.610 0.433 ;
      RECT 0.217 0.698 0.610 0.812 ;
      RECT 0.242 0.294 0.589 0.408 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.150 0.487 0.376 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.557 -0.080 1.100 0.080 ;
      RECT 0.463 -0.080 0.557 0.218 ;
      RECT 0.156 -0.080 0.463 0.080 ;
      RECT 0.061 -0.080 0.156 0.122 ;
      RECT 0.000 -0.080 0.061 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.922 1.120 1.100 1.280 ;
      RECT 0.828 0.917 0.922 1.280 ;
      RECT 0.532 1.120 0.828 1.280 ;
      RECT 0.438 0.917 0.532 1.280 ;
      RECT 0.144 1.120 0.438 1.280 ;
      RECT 0.050 0.917 0.144 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
END CLKINVX8

MACRO CLKINVX4
  CLASS CORE ;
  FOREIGN CLKINVX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.307 0.488 0.900 ;
      RECT 0.286 0.307 0.387 0.398 ;
      RECT 0.382 0.706 0.387 0.900 ;
      RECT 0.292 0.706 0.382 1.001 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.481 0.252 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.647 -0.080 0.700 0.080 ;
      RECT 0.557 -0.080 0.647 0.122 ;
      RECT 0.180 -0.080 0.557 0.080 ;
      RECT 0.090 -0.080 0.180 0.122 ;
      RECT 0.000 -0.080 0.090 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.583 1.120 0.700 1.280 ;
      RECT 0.493 1.078 0.583 1.280 ;
      RECT 0.180 1.120 0.493 1.280 ;
      RECT 0.090 1.078 0.180 1.280 ;
      RECT 0.000 1.120 0.090 1.280 ;
     END
  END VDD
END CLKINVX4

MACRO CLKINVX3
  CLASS CORE ;
  FOREIGN CLKINVX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.311 0.626 0.358 0.900 ;
      RECT 0.241 0.342 0.311 0.900 ;
      RECT 0.223 0.627 0.241 0.900 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.162 0.581 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.497 -0.080 0.600 0.080 ;
      RECT 0.394 -0.080 0.497 0.122 ;
      RECT 0.000 -0.080 0.394 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.158 1.120 0.600 1.280 ;
      RECT 0.055 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.055 1.280 ;
     END
  END VDD
END CLKINVX3

MACRO CLKINVX2
  CLASS CORE ;
  FOREIGN CLKINVX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.400 0.286 0.470 0.787 ;
      RECT 0.350 0.286 0.400 0.367 ;
      RECT 0.224 0.700 0.400 0.787 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.329 0.574 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.220 -0.080 0.600 0.080 ;
      RECT 0.117 -0.080 0.220 0.352 ;
      RECT 0.000 -0.080 0.117 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.439 1.120 0.600 1.280 ;
      RECT 0.324 1.061 0.439 1.280 ;
      RECT 0.000 1.120 0.324 1.280 ;
     END
  END VDD
END CLKINVX2

MACRO CLKINVX20
  CLASS CORE ;
  FOREIGN CLKINVX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.867 0.696 5.033 0.889 ;
      RECT 4.454 0.286 4.867 0.900 ;
      RECT 2.371 0.285 4.454 0.436 ;
      RECT 4.278 0.712 4.454 0.874 ;
      RECT 4.127 0.696 4.278 0.889 ;
      RECT 3.926 0.712 4.127 0.874 ;
      RECT 3.762 0.696 3.926 0.889 ;
      RECT 3.479 0.712 3.762 0.874 ;
      RECT 3.388 0.696 3.479 0.889 ;
      RECT 3.096 0.712 3.388 0.874 ;
      RECT 2.932 0.696 3.096 0.889 ;
      RECT 2.718 0.712 2.932 0.874 ;
      RECT 2.581 0.696 2.718 0.889 ;
      RECT 2.343 0.712 2.581 0.874 ;
      RECT 2.229 0.696 2.343 0.889 ;
      RECT 1.992 0.712 2.229 0.874 ;
      RECT 1.868 0.696 1.992 0.889 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.191 0.500 0.314 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.205 -0.080 5.100 0.080 ;
      RECT 4.114 -0.080 4.205 0.214 ;
      RECT 3.836 -0.080 4.114 0.080 ;
      RECT 3.745 -0.080 3.836 0.214 ;
      RECT 3.457 -0.080 3.745 0.080 ;
      RECT 3.367 -0.080 3.457 0.214 ;
      RECT 3.076 -0.080 3.367 0.080 ;
      RECT 2.986 -0.080 3.076 0.214 ;
      RECT 2.698 -0.080 2.986 0.080 ;
      RECT 2.607 -0.080 2.698 0.214 ;
      RECT 2.320 -0.080 2.607 0.080 ;
      RECT 2.229 -0.080 2.320 0.214 ;
      RECT 1.382 -0.080 2.229 0.080 ;
      RECT 1.291 -0.080 1.382 0.210 ;
      RECT 0.970 -0.080 1.291 0.080 ;
      RECT 0.879 -0.080 0.970 0.210 ;
      RECT 0.590 -0.080 0.879 0.080 ;
      RECT 0.500 -0.080 0.590 0.223 ;
      RECT 0.000 -0.080 0.500 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.800 1.120 5.100 1.280 ;
      RECT 4.710 0.996 4.800 1.280 ;
      RECT 4.421 1.120 4.710 1.280 ;
      RECT 4.330 0.996 4.421 1.280 ;
      RECT 4.042 1.120 4.330 1.280 ;
      RECT 3.952 0.996 4.042 1.280 ;
      RECT 3.662 1.120 3.952 1.280 ;
      RECT 3.572 0.996 3.662 1.280 ;
      RECT 3.287 1.120 3.572 1.280 ;
      RECT 3.196 0.996 3.287 1.280 ;
      RECT 2.908 1.120 3.196 1.280 ;
      RECT 2.818 0.983 2.908 1.280 ;
      RECT 2.526 1.120 2.818 1.280 ;
      RECT 2.435 0.983 2.526 1.280 ;
      RECT 2.148 1.120 2.435 1.280 ;
      RECT 2.057 0.983 2.148 1.280 ;
      RECT 1.769 1.120 2.057 1.280 ;
      RECT 1.679 0.985 1.769 1.280 ;
      RECT 1.351 1.120 1.679 1.280 ;
      RECT 1.260 0.982 1.351 1.280 ;
      RECT 0.969 1.120 1.260 1.280 ;
      RECT 0.878 0.982 0.969 1.280 ;
      RECT 0.577 1.120 0.878 1.280 ;
      RECT 0.486 0.989 0.577 1.280 ;
      RECT 0.214 1.120 0.486 1.280 ;
      RECT 0.124 0.741 0.214 1.280 ;
      RECT 0.000 1.120 0.124 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.691 0.505 4.318 0.640 ;
      RECT 1.547 0.281 1.691 0.821 ;
      RECT 1.519 0.281 1.547 0.875 ;
      RECT 0.690 0.281 1.519 0.435 ;
      RECT 1.456 0.668 1.519 0.875 ;
      RECT 1.158 0.668 1.456 0.821 ;
      RECT 0.630 0.500 1.347 0.581 ;
      RECT 1.067 0.668 1.158 0.889 ;
      RECT 0.779 0.668 1.067 0.821 ;
      RECT 0.690 0.668 0.779 0.889 ;
      RECT 0.689 0.696 0.690 0.889 ;
      RECT 0.437 0.513 0.630 0.568 ;
      RECT 0.376 0.343 0.437 0.789 ;
      RECT 0.326 0.343 0.376 0.424 ;
      RECT 0.329 0.708 0.376 0.789 ;
  END
END CLKINVX20

MACRO CLKINVX16
  CLASS CORE ;
  FOREIGN CLKINVX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.929 0.286 4.343 0.914 ;
      RECT 3.464 0.286 3.929 0.448 ;
      RECT 3.785 0.712 3.929 0.874 ;
      RECT 3.639 0.696 3.785 0.889 ;
      RECT 3.411 0.712 3.639 0.874 ;
      RECT 3.121 0.285 3.464 0.448 ;
      RECT 3.287 0.696 3.411 0.889 ;
      RECT 3.049 0.712 3.287 0.874 ;
      RECT 2.185 0.286 3.121 0.448 ;
      RECT 2.935 0.696 3.049 0.889 ;
      RECT 2.697 0.712 2.935 0.874 ;
      RECT 2.559 0.696 2.697 0.889 ;
      RECT 2.345 0.712 2.559 0.874 ;
      RECT 2.177 0.696 2.345 0.889 ;
      RECT 1.889 0.712 2.177 0.874 ;
      RECT 1.799 0.696 1.889 0.889 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.191 0.500 0.315 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.641 -0.080 4.400 0.080 ;
      RECT 3.551 -0.080 3.641 0.214 ;
      RECT 3.272 -0.080 3.551 0.080 ;
      RECT 3.181 -0.080 3.272 0.214 ;
      RECT 2.893 -0.080 3.181 0.080 ;
      RECT 2.803 -0.080 2.893 0.214 ;
      RECT 2.512 -0.080 2.803 0.080 ;
      RECT 2.421 -0.080 2.512 0.214 ;
      RECT 2.133 -0.080 2.421 0.080 ;
      RECT 2.043 -0.080 2.133 0.214 ;
      RECT 0.971 -0.080 2.043 0.080 ;
      RECT 0.880 -0.080 0.971 0.228 ;
      RECT 0.591 -0.080 0.880 0.080 ;
      RECT 0.500 -0.080 0.591 0.223 ;
      RECT 0.000 -0.080 0.500 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.331 1.120 4.400 1.280 ;
      RECT 4.240 0.996 4.331 1.280 ;
      RECT 3.975 1.120 4.240 1.280 ;
      RECT 3.884 0.996 3.975 1.280 ;
      RECT 3.595 1.120 3.884 1.280 ;
      RECT 3.504 0.996 3.595 1.280 ;
      RECT 3.219 1.120 3.504 1.280 ;
      RECT 3.128 0.996 3.219 1.280 ;
      RECT 2.840 1.120 3.128 1.280 ;
      RECT 2.749 0.983 2.840 1.280 ;
      RECT 2.457 1.120 2.749 1.280 ;
      RECT 2.367 0.983 2.457 1.280 ;
      RECT 2.079 1.120 2.367 1.280 ;
      RECT 1.988 0.983 2.079 1.280 ;
      RECT 1.700 1.120 1.988 1.280 ;
      RECT 1.609 0.985 1.700 1.280 ;
      RECT 1.352 1.120 1.609 1.280 ;
      RECT 1.261 0.982 1.352 1.280 ;
      RECT 0.969 1.120 1.261 1.280 ;
      RECT 0.879 0.982 0.969 1.280 ;
      RECT 0.577 1.120 0.879 1.280 ;
      RECT 0.487 0.989 0.577 1.280 ;
      RECT 0.215 1.120 0.487 1.280 ;
      RECT 0.124 0.741 0.215 1.280 ;
      RECT 0.000 1.120 0.124 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.717 0.521 3.813 0.602 ;
      RECT 1.605 0.526 1.717 0.598 ;
      RECT 1.424 0.319 1.605 0.807 ;
      RECT 0.689 0.319 1.424 0.445 ;
      RECT 1.159 0.643 1.424 0.807 ;
      RECT 0.607 0.500 1.324 0.581 ;
      RECT 1.068 0.643 1.159 0.889 ;
      RECT 0.780 0.643 1.068 0.807 ;
      RECT 0.689 0.643 0.780 0.889 ;
      RECT 0.437 0.513 0.607 0.568 ;
      RECT 0.376 0.343 0.437 0.789 ;
      RECT 0.327 0.343 0.376 0.424 ;
      RECT 0.329 0.708 0.376 0.789 ;
  END
END CLKINVX16

MACRO CLKBUFXL
  CLASS CORE ;
  FOREIGN CLKBUFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.582 0.290 0.643 0.712 ;
      RECT 0.509 0.290 0.582 0.345 ;
      RECT 0.562 0.627 0.582 0.712 ;
      RECT 0.498 0.657 0.562 0.712 ;
      RECT 0.419 0.264 0.509 0.345 ;
      RECT 0.408 0.657 0.498 0.738 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.215 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.323 1.120 0.700 1.280 ;
      RECT 0.233 1.078 0.323 1.280 ;
      RECT 0.000 1.120 0.233 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.337 0.433 0.403 0.514 ;
      RECT 0.276 0.290 0.337 0.712 ;
      RECT 0.138 0.290 0.276 0.345 ;
      RECT 0.138 0.657 0.276 0.712 ;
      RECT 0.048 0.264 0.138 0.345 ;
      RECT 0.048 0.657 0.138 0.738 ;
  END
END CLKBUFXL

MACRO CLKBUFX8
  CLASS CORE ;
  FOREIGN CLKBUFX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.126 0.433 1.240 0.767 ;
      RECT 0.803 0.321 1.126 0.767 ;
      RECT 0.782 0.321 0.803 0.440 ;
      RECT 0.782 0.625 0.803 0.757 ;
      RECT 0.636 0.321 0.782 0.402 ;
      RECT 0.613 0.676 0.782 0.757 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.311 0.474 0.391 0.555 ;
      RECT 0.246 0.439 0.311 0.555 ;
      RECT 0.160 0.474 0.246 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.912 -0.080 1.300 0.080 ;
      RECT 0.816 -0.080 0.912 0.215 ;
      RECT 0.552 -0.080 0.816 0.080 ;
      RECT 0.456 -0.080 0.552 0.215 ;
      RECT 0.000 -0.080 0.456 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 1.120 1.300 1.280 ;
      RECT 1.154 0.877 1.249 1.280 ;
      RECT 0.889 1.120 1.154 1.280 ;
      RECT 0.794 0.877 0.889 1.280 ;
      RECT 0.518 1.120 0.794 1.280 ;
      RECT 0.422 1.078 0.518 1.280 ;
      RECT 0.146 1.120 0.422 1.280 ;
      RECT 0.051 0.844 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.549 0.519 0.718 0.600 ;
      RECT 0.484 0.300 0.549 0.712 ;
      RECT 0.349 0.300 0.484 0.355 ;
      RECT 0.326 0.657 0.484 0.712 ;
      RECT 0.253 0.274 0.349 0.355 ;
      RECT 0.231 0.657 0.326 0.738 ;
  END
END CLKBUFX8

MACRO CLKBUFX4
  CLASS CORE ;
  FOREIGN CLKBUFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.641 0.300 0.682 0.633 ;
      RECT 0.578 0.300 0.641 0.714 ;
      RECT 0.464 0.331 0.578 0.412 ;
      RECT 0.556 0.660 0.578 0.714 ;
      RECT 0.464 0.660 0.556 0.740 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.433 0.221 0.570 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.764 -0.080 0.900 0.080 ;
      RECT 0.671 -0.080 0.764 0.122 ;
      RECT 0.322 -0.080 0.671 0.080 ;
      RECT 0.229 -0.080 0.322 0.122 ;
      RECT 0.000 -0.080 0.229 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.764 1.120 0.900 1.280 ;
      RECT 0.671 1.078 0.764 1.280 ;
      RECT 0.349 1.120 0.671 1.280 ;
      RECT 0.334 1.078 0.349 1.280 ;
      RECT 0.271 1.065 0.334 1.280 ;
      RECT 0.256 1.078 0.271 1.280 ;
      RECT 0.000 1.120 0.256 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.346 0.490 0.515 0.571 ;
      RECT 0.284 0.324 0.346 0.707 ;
      RECT 0.142 0.324 0.284 0.379 ;
      RECT 0.142 0.652 0.284 0.707 ;
      RECT 0.049 0.298 0.142 0.379 ;
      RECT 0.049 0.652 0.142 0.733 ;
  END
END CLKBUFX4

MACRO CLKBUFX3
  CLASS CORE ;
  FOREIGN CLKBUFX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.469 0.287 0.498 0.368 ;
      RECT 0.469 0.433 0.488 0.752 ;
      RECT 0.408 0.287 0.469 0.752 ;
      RECT 0.398 0.433 0.408 0.752 ;
      RECT 0.387 0.433 0.398 0.633 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.433 0.147 0.562 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 -0.080 0.700 0.080 ;
      RECT 0.562 -0.080 0.652 0.122 ;
      RECT 0.313 -0.080 0.562 0.080 ;
      RECT 0.223 -0.080 0.313 0.122 ;
      RECT 0.000 -0.080 0.223 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 1.120 0.700 1.280 ;
      RECT 0.562 1.078 0.652 1.280 ;
      RECT 0.317 1.120 0.562 1.280 ;
      RECT 0.215 1.078 0.317 1.280 ;
      RECT 0.000 1.120 0.215 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.296 0.470 0.325 0.551 ;
      RECT 0.235 0.270 0.296 0.751 ;
      RECT 0.138 0.270 0.235 0.325 ;
      RECT 0.138 0.696 0.235 0.751 ;
      RECT 0.048 0.244 0.138 0.325 ;
      RECT 0.048 0.696 0.138 0.777 ;
  END
END CLKBUFX3

MACRO CLKBUFX2
  CLASS CORE ;
  FOREIGN CLKBUFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.583 0.301 0.643 0.710 ;
      RECT 0.582 0.275 0.583 0.710 ;
      RECT 0.435 0.275 0.582 0.356 ;
      RECT 0.562 0.627 0.582 0.736 ;
      RECT 0.424 0.655 0.562 0.736 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.239 0.538 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.323 -0.080 0.700 0.080 ;
      RECT 0.233 -0.080 0.323 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.298 1.078 0.313 1.280 ;
      RECT 0.237 1.065 0.298 1.280 ;
      RECT 0.223 1.078 0.237 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.363 0.490 0.430 0.571 ;
      RECT 0.302 0.301 0.363 0.710 ;
      RECT 0.164 0.301 0.302 0.356 ;
      RECT 0.164 0.655 0.302 0.710 ;
      RECT 0.074 0.275 0.164 0.356 ;
      RECT 0.074 0.655 0.164 0.736 ;
  END
END CLKBUFX2

MACRO CLKBUFX20
  CLASS CORE ;
  FOREIGN CLKBUFX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.914 0.286 3.968 0.914 ;
      RECT 3.557 0.268 3.914 0.914 ;
      RECT 1.246 0.268 3.557 0.448 ;
      RECT 3.537 0.633 3.557 0.839 ;
      RECT 1.236 0.659 3.537 0.839 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.818 0.474 0.992 0.555 ;
      RECT 0.757 0.439 0.818 0.555 ;
      RECT 0.154 0.474 0.757 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.864 -0.080 4.200 0.080 ;
      RECT 2.773 -0.080 2.864 0.198 ;
      RECT 2.524 -0.080 2.773 0.080 ;
      RECT 2.434 -0.080 2.524 0.198 ;
      RECT 2.185 -0.080 2.434 0.080 ;
      RECT 2.095 -0.080 2.185 0.198 ;
      RECT 1.845 -0.080 2.095 0.080 ;
      RECT 1.755 -0.080 1.845 0.198 ;
      RECT 1.506 -0.080 1.755 0.080 ;
      RECT 1.416 -0.080 1.506 0.198 ;
      RECT 1.167 -0.080 1.416 0.080 ;
      RECT 1.077 -0.080 1.167 0.214 ;
      RECT 0.785 -0.080 1.077 0.080 ;
      RECT 0.695 -0.080 0.785 0.214 ;
      RECT 0.403 -0.080 0.695 0.080 ;
      RECT 0.313 -0.080 0.403 0.214 ;
      RECT 0.000 -0.080 0.313 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.882 1.120 4.200 1.280 ;
      RECT 3.867 1.078 3.882 1.280 ;
      RECT 3.806 1.065 3.867 1.280 ;
      RECT 3.792 1.078 3.806 1.280 ;
      RECT 3.532 1.120 3.792 1.280 ;
      RECT 3.442 0.989 3.532 1.280 ;
      RECT 3.192 1.120 3.442 1.280 ;
      RECT 3.102 0.989 3.192 1.280 ;
      RECT 2.853 1.120 3.102 1.280 ;
      RECT 2.763 0.989 2.853 1.280 ;
      RECT 2.514 1.120 2.763 1.280 ;
      RECT 2.423 0.989 2.514 1.280 ;
      RECT 2.174 1.120 2.423 1.280 ;
      RECT 2.084 0.989 2.174 1.280 ;
      RECT 1.835 1.120 2.084 1.280 ;
      RECT 1.745 0.972 1.835 1.280 ;
      RECT 1.495 1.120 1.745 1.280 ;
      RECT 1.405 0.972 1.495 1.280 ;
      RECT 1.156 1.120 1.405 1.280 ;
      RECT 1.066 0.954 1.156 1.280 ;
      RECT 0.817 1.120 1.066 1.280 ;
      RECT 0.727 0.954 0.817 1.280 ;
      RECT 0.477 1.120 0.727 1.280 ;
      RECT 0.387 0.954 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.954 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.172 0.513 3.426 0.594 ;
      RECT 1.082 0.283 1.172 0.757 ;
      RECT 0.504 0.283 1.082 0.364 ;
      RECT 0.217 0.676 1.082 0.757 ;
  END
END CLKBUFX20

MACRO CLKBUFX1
  CLASS CORE ;
  FOREIGN CLKBUFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.582 0.290 0.643 0.726 ;
      RECT 0.509 0.290 0.582 0.345 ;
      RECT 0.562 0.627 0.582 0.726 ;
      RECT 0.488 0.671 0.562 0.726 ;
      RECT 0.419 0.264 0.509 0.345 ;
      RECT 0.398 0.671 0.488 0.752 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.215 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.223 1.078 0.313 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.337 0.490 0.403 0.571 ;
      RECT 0.276 0.290 0.337 0.712 ;
      RECT 0.138 0.290 0.276 0.345 ;
      RECT 0.138 0.657 0.276 0.712 ;
      RECT 0.048 0.264 0.138 0.345 ;
      RECT 0.048 0.657 0.138 0.738 ;
  END
END CLKBUFX1

MACRO CLKBUFX16
  CLASS CORE ;
  FOREIGN CLKBUFX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.189 0.286 3.243 0.914 ;
      RECT 2.836 0.268 3.189 0.914 ;
      RECT 1.068 0.268 2.836 0.448 ;
      RECT 2.816 0.633 2.836 0.839 ;
      RECT 1.084 0.659 2.816 0.839 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.337 0.426 0.797 0.507 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.389 -0.080 3.300 0.080 ;
      RECT 2.300 -0.080 2.389 0.198 ;
      RECT 2.011 -0.080 2.300 0.080 ;
      RECT 1.921 -0.080 2.011 0.198 ;
      RECT 1.663 -0.080 1.921 0.080 ;
      RECT 1.574 -0.080 1.663 0.198 ;
      RECT 1.326 -0.080 1.574 0.080 ;
      RECT 1.237 -0.080 1.326 0.198 ;
      RECT 0.989 -0.080 1.237 0.080 ;
      RECT 0.900 -0.080 0.989 0.198 ;
      RECT 0.611 -0.080 0.900 0.080 ;
      RECT 0.521 -0.080 0.611 0.198 ;
      RECT 0.000 -0.080 0.521 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.047 1.120 3.300 1.280 ;
      RECT 2.958 0.989 3.047 1.280 ;
      RECT 2.700 1.120 2.958 1.280 ;
      RECT 2.611 0.972 2.700 1.280 ;
      RECT 2.363 1.120 2.611 1.280 ;
      RECT 2.274 0.972 2.363 1.280 ;
      RECT 2.026 1.120 2.274 1.280 ;
      RECT 1.937 0.972 2.026 1.280 ;
      RECT 1.679 1.120 1.937 1.280 ;
      RECT 1.589 0.972 1.679 1.280 ;
      RECT 1.342 1.120 1.589 1.280 ;
      RECT 1.253 0.972 1.342 1.280 ;
      RECT 1.005 1.120 1.253 1.280 ;
      RECT 0.916 0.972 1.005 1.280 ;
      RECT 0.658 1.120 0.916 1.280 ;
      RECT 0.568 0.877 0.658 1.280 ;
      RECT 0.311 1.120 0.568 1.280 ;
      RECT 0.296 1.078 0.311 1.280 ;
      RECT 0.236 1.065 0.296 1.280 ;
      RECT 0.221 1.078 0.236 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.995 0.513 2.726 0.594 ;
      RECT 0.905 0.274 0.995 0.738 ;
      RECT 0.332 0.274 0.905 0.355 ;
      RECT 0.400 0.657 0.905 0.738 ;
  END
END CLKBUFX16

MACRO BUFXL
  CLASS CORE ;
  FOREIGN BUFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.582 0.274 0.643 0.726 ;
      RECT 0.498 0.274 0.582 0.329 ;
      RECT 0.562 0.627 0.582 0.726 ;
      RECT 0.488 0.671 0.562 0.726 ;
      RECT 0.408 0.248 0.498 0.329 ;
      RECT 0.398 0.671 0.488 0.752 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.215 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.223 1.078 0.313 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.337 0.490 0.403 0.571 ;
      RECT 0.276 0.290 0.337 0.712 ;
      RECT 0.138 0.290 0.276 0.345 ;
      RECT 0.138 0.657 0.276 0.712 ;
      RECT 0.048 0.264 0.138 0.345 ;
      RECT 0.048 0.657 0.138 0.738 ;
  END
END BUFXL

MACRO BUFX8
  CLASS CORE ;
  FOREIGN BUFX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.220 0.433 1.364 0.767 ;
      RECT 1.131 0.433 1.220 0.774 ;
      RECT 0.947 0.307 1.131 0.774 ;
      RECT 0.927 0.307 0.947 0.440 ;
      RECT 0.927 0.626 0.947 0.774 ;
      RECT 0.609 0.307 0.927 0.421 ;
      RECT 0.587 0.660 0.927 0.774 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.298 0.474 0.372 0.555 ;
      RECT 0.236 0.439 0.298 0.555 ;
      RECT 0.154 0.474 0.236 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.218 -0.080 1.600 0.080 ;
      RECT 1.126 -0.080 1.218 0.211 ;
      RECT 0.873 -0.080 1.126 0.080 ;
      RECT 0.781 -0.080 0.873 0.211 ;
      RECT 0.528 -0.080 0.781 0.080 ;
      RECT 0.436 -0.080 0.528 0.198 ;
      RECT 0.140 -0.080 0.436 0.080 ;
      RECT 0.048 -0.080 0.140 0.211 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.196 1.120 1.600 1.280 ;
      RECT 1.104 0.877 1.196 1.280 ;
      RECT 0.851 1.120 1.104 1.280 ;
      RECT 0.760 0.877 0.851 1.280 ;
      RECT 0.506 1.120 0.760 1.280 ;
      RECT 0.415 0.897 0.506 1.280 ;
      RECT 0.162 1.120 0.415 1.280 ;
      RECT 0.070 0.897 0.162 1.280 ;
      RECT 0.000 1.120 0.070 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.525 0.519 0.865 0.600 ;
      RECT 0.434 0.274 0.525 0.738 ;
      RECT 0.242 0.274 0.434 0.355 ;
      RECT 0.242 0.657 0.434 0.738 ;
  END
END BUFX8

MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.600 0.300 0.682 0.733 ;
      RECT 0.578 0.300 0.600 0.767 ;
      RECT 0.556 0.300 0.578 0.412 ;
      RECT 0.556 0.652 0.578 0.767 ;
      RECT 0.464 0.219 0.556 0.412 ;
      RECT 0.464 0.652 0.556 0.957 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.433 0.218 0.570 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.764 -0.080 0.900 0.080 ;
      RECT 0.671 -0.080 0.764 0.122 ;
      RECT 0.349 -0.080 0.671 0.080 ;
      RECT 0.256 -0.080 0.349 0.122 ;
      RECT 0.000 -0.080 0.256 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.764 1.120 0.900 1.280 ;
      RECT 0.671 0.953 0.764 1.280 ;
      RECT 0.349 1.120 0.671 1.280 ;
      RECT 0.256 0.953 0.349 1.280 ;
      RECT 0.000 1.120 0.256 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.376 0.477 0.515 0.585 ;
      RECT 0.284 0.298 0.376 0.733 ;
      RECT 0.142 0.298 0.284 0.379 ;
      RECT 0.142 0.652 0.284 0.733 ;
      RECT 0.049 0.186 0.142 0.379 ;
      RECT 0.049 0.652 0.142 0.957 ;
  END
END BUFX4

MACRO BUFX3
  CLASS CORE ;
  FOREIGN BUFX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.469 0.287 0.498 0.368 ;
      RECT 0.469 0.433 0.488 0.752 ;
      RECT 0.408 0.287 0.469 0.752 ;
      RECT 0.398 0.433 0.408 0.752 ;
      RECT 0.387 0.433 0.398 0.633 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.433 0.147 0.562 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.647 -0.080 0.700 0.080 ;
      RECT 0.557 -0.080 0.647 0.122 ;
      RECT 0.000 -0.080 0.557 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.286 1.120 0.700 1.280 ;
      RECT 0.196 1.078 0.286 1.280 ;
      RECT 0.000 1.120 0.196 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.296 0.470 0.325 0.551 ;
      RECT 0.235 0.270 0.296 0.751 ;
      RECT 0.138 0.270 0.235 0.325 ;
      RECT 0.138 0.696 0.235 0.751 ;
      RECT 0.048 0.244 0.138 0.325 ;
      RECT 0.048 0.696 0.138 0.777 ;
  END
END BUFX3

MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.623 0.439 0.643 0.494 ;
      RECT 0.562 0.357 0.623 0.710 ;
      RECT 0.525 0.357 0.562 0.412 ;
      RECT 0.514 0.655 0.562 0.710 ;
      RECT 0.435 0.331 0.525 0.412 ;
      RECT 0.424 0.655 0.514 0.736 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.236 0.538 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.323 -0.080 0.700 0.080 ;
      RECT 0.233 -0.080 0.323 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.298 1.078 0.313 1.280 ;
      RECT 0.237 1.065 0.298 1.280 ;
      RECT 0.223 1.078 0.237 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.363 0.490 0.430 0.571 ;
      RECT 0.302 0.301 0.363 0.712 ;
      RECT 0.164 0.301 0.302 0.356 ;
      RECT 0.164 0.657 0.302 0.712 ;
      RECT 0.074 0.275 0.164 0.356 ;
      RECT 0.074 0.657 0.164 0.738 ;
  END
END BUFX2

MACRO BUFX20
  CLASS CORE ;
  FOREIGN BUFX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.332 0.268 2.743 0.914 ;
      RECT 0.907 0.268 2.332 0.408 ;
      RECT 2.312 0.683 2.332 0.839 ;
      RECT 0.896 0.699 2.312 0.839 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.468 0.474 0.663 0.555 ;
      RECT 0.407 0.439 0.468 0.555 ;
      RECT 0.199 0.474 0.407 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.535 -0.080 2.800 0.080 ;
      RECT 2.445 -0.080 2.535 0.122 ;
      RECT 2.185 -0.080 2.445 0.080 ;
      RECT 2.095 -0.080 2.185 0.198 ;
      RECT 1.845 -0.080 2.095 0.080 ;
      RECT 1.755 -0.080 1.845 0.198 ;
      RECT 1.506 -0.080 1.755 0.080 ;
      RECT 1.416 -0.080 1.506 0.198 ;
      RECT 1.167 -0.080 1.416 0.080 ;
      RECT 1.077 -0.080 1.167 0.198 ;
      RECT 0.827 -0.080 1.077 0.080 ;
      RECT 0.737 -0.080 0.827 0.215 ;
      RECT 0.477 -0.080 0.737 0.080 ;
      RECT 0.387 -0.080 0.477 0.234 ;
      RECT 0.138 -0.080 0.387 0.080 ;
      RECT 0.048 -0.080 0.138 0.234 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.524 1.120 2.800 1.280 ;
      RECT 2.510 1.078 2.524 1.280 ;
      RECT 2.449 1.065 2.510 1.280 ;
      RECT 2.434 1.078 2.449 1.280 ;
      RECT 2.174 1.120 2.434 1.280 ;
      RECT 2.084 0.989 2.174 1.280 ;
      RECT 1.835 1.120 2.084 1.280 ;
      RECT 1.745 0.989 1.835 1.280 ;
      RECT 1.495 1.120 1.745 1.280 ;
      RECT 1.405 0.972 1.495 1.280 ;
      RECT 1.156 1.120 1.405 1.280 ;
      RECT 1.066 0.972 1.156 1.280 ;
      RECT 0.817 1.120 1.066 1.280 ;
      RECT 0.727 0.873 0.817 1.280 ;
      RECT 0.477 1.120 0.727 1.280 ;
      RECT 0.387 0.873 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.873 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.834 0.513 2.190 0.594 ;
      RECT 0.744 0.320 0.834 0.757 ;
      RECT 0.557 0.320 0.744 0.401 ;
      RECT 0.217 0.676 0.744 0.757 ;
      RECT 0.308 0.320 0.557 0.375 ;
      RECT 0.217 0.320 0.308 0.401 ;
  END
END BUFX20

MACRO BUFX1
  CLASS CORE ;
  FOREIGN BUFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.582 0.274 0.643 0.726 ;
      RECT 0.498 0.274 0.582 0.329 ;
      RECT 0.562 0.627 0.582 0.726 ;
      RECT 0.488 0.671 0.562 0.726 ;
      RECT 0.408 0.248 0.498 0.329 ;
      RECT 0.398 0.671 0.488 0.752 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.215 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.297 -0.080 0.700 0.080 ;
      RECT 0.207 -0.080 0.297 0.122 ;
      RECT 0.000 -0.080 0.207 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.223 1.078 0.313 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.337 0.490 0.403 0.571 ;
      RECT 0.276 0.290 0.337 0.712 ;
      RECT 0.138 0.290 0.276 0.345 ;
      RECT 0.138 0.657 0.276 0.712 ;
      RECT 0.048 0.264 0.138 0.345 ;
      RECT 0.048 0.657 0.138 0.738 ;
  END
END BUFX1

MACRO BUFX16
  CLASS CORE ;
  FOREIGN BUFX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.827 0.268 2.242 0.914 ;
      RECT 0.745 0.268 1.827 0.408 ;
      RECT 1.807 0.675 1.827 0.839 ;
      RECT 0.917 0.699 1.807 0.839 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.473 0.521 0.547 0.602 ;
      RECT 0.411 0.521 0.473 0.627 ;
      RECT 0.155 0.521 0.411 0.602 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.069 -0.080 2.300 0.080 ;
      RECT 1.978 -0.080 2.069 0.122 ;
      RECT 1.705 -0.080 1.978 0.080 ;
      RECT 1.614 -0.080 1.705 0.198 ;
      RECT 1.351 -0.080 1.614 0.080 ;
      RECT 1.260 -0.080 1.351 0.198 ;
      RECT 1.008 -0.080 1.260 0.080 ;
      RECT 0.917 -0.080 1.008 0.198 ;
      RECT 0.654 -0.080 0.917 0.080 ;
      RECT 0.563 -0.080 0.654 0.216 ;
      RECT 0.311 -0.080 0.563 0.080 ;
      RECT 0.220 -0.080 0.311 0.215 ;
      RECT 0.000 -0.080 0.220 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.252 1.120 2.300 1.280 ;
      RECT 2.161 1.078 2.252 1.280 ;
      RECT 1.887 1.120 2.161 1.280 ;
      RECT 1.796 1.078 1.887 1.280 ;
      RECT 1.523 1.120 1.796 1.280 ;
      RECT 1.431 0.972 1.523 1.280 ;
      RECT 1.179 1.120 1.431 1.280 ;
      RECT 1.088 0.972 1.179 1.280 ;
      RECT 0.836 1.120 1.088 1.280 ;
      RECT 0.745 0.972 0.836 1.280 ;
      RECT 0.483 1.120 0.745 1.280 ;
      RECT 0.391 0.823 0.483 1.280 ;
      RECT 0.139 1.120 0.391 1.280 ;
      RECT 0.048 0.823 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.672 0.513 1.745 0.594 ;
      RECT 0.610 0.335 0.672 0.743 ;
      RECT 0.048 0.335 0.610 0.415 ;
      RECT 0.563 0.657 0.610 0.743 ;
      RECT 0.311 0.688 0.563 0.743 ;
      RECT 0.220 0.657 0.311 0.743 ;
  END
END BUFX16

MACRO BUFX12
  CLASS CORE ;
  FOREIGN BUFX12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.319 0.300 1.741 0.767 ;
      RECT 1.298 0.321 1.319 0.440 ;
      RECT 1.298 0.626 1.319 0.757 ;
      RECT 0.769 0.321 1.298 0.402 ;
      RECT 0.747 0.676 1.298 0.757 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.301 0.474 0.554 0.555 ;
      RECT 0.239 0.439 0.301 0.555 ;
      RECT 0.194 0.474 0.239 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.735 -0.080 1.800 0.080 ;
      RECT 1.642 -0.080 1.735 0.211 ;
      RECT 1.385 -0.080 1.642 0.080 ;
      RECT 1.293 -0.080 1.385 0.211 ;
      RECT 1.036 -0.080 1.293 0.080 ;
      RECT 0.944 -0.080 1.036 0.215 ;
      RECT 0.687 -0.080 0.944 0.080 ;
      RECT 0.595 -0.080 0.687 0.215 ;
      RECT 0.327 -0.080 0.595 0.080 ;
      RECT 0.235 -0.080 0.327 0.122 ;
      RECT 0.000 -0.080 0.235 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.751 1.120 1.800 1.280 ;
      RECT 1.658 0.972 1.751 1.280 ;
      RECT 1.377 1.120 1.658 1.280 ;
      RECT 1.285 0.972 1.377 1.280 ;
      RECT 1.015 1.120 1.285 1.280 ;
      RECT 0.922 0.972 1.015 1.280 ;
      RECT 0.665 1.120 0.922 1.280 ;
      RECT 0.573 0.897 0.665 1.280 ;
      RECT 0.316 1.120 0.573 1.280 ;
      RECT 0.224 0.897 0.316 1.280 ;
      RECT 0.000 1.120 0.224 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.685 0.519 1.193 0.600 ;
      RECT 0.622 0.345 0.685 0.712 ;
      RECT 0.513 0.345 0.622 0.400 ;
      RECT 0.491 0.657 0.622 0.712 ;
      RECT 0.420 0.319 0.513 0.400 ;
      RECT 0.398 0.657 0.491 0.738 ;
      RECT 0.142 0.319 0.420 0.374 ;
      RECT 0.142 0.657 0.398 0.712 ;
      RECT 0.079 0.319 0.142 0.389 ;
      RECT 0.049 0.657 0.142 0.738 ;
      RECT 0.049 0.335 0.079 0.389 ;
  END
END BUFX12

MACRO AOI33X1
  CLASS CORE ;
  FOREIGN AOI33X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.323 0.573 1.343 0.627 ;
      RECT 1.282 0.215 1.323 0.746 ;
      RECT 1.262 0.215 1.282 0.767 ;
      RECT 0.536 0.215 1.262 0.270 ;
      RECT 1.252 0.692 1.262 0.767 ;
      RECT 1.161 0.692 1.252 0.912 ;
      RECT 0.932 0.692 1.161 0.746 ;
      RECT 0.780 0.692 0.932 0.773 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.419 0.223 0.511 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.199 0.567 0.391 0.660 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.377 0.395 0.566 0.500 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.034 0.383 1.168 0.507 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.933 0.567 1.038 0.633 ;
      RECT 0.843 0.546 0.933 0.633 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.639 0.546 0.776 0.633 ;
      RECT 0.582 0.573 0.639 0.627 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.124 -0.080 1.400 0.080 ;
      RECT 1.034 -0.080 1.124 0.122 ;
      RECT 0.138 -0.080 1.034 0.080 ;
      RECT 0.048 -0.080 0.138 0.325 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.530 1.120 1.400 1.280 ;
      RECT 0.440 1.078 0.530 1.280 ;
      RECT 0.138 1.120 0.440 1.280 ;
      RECT 0.048 0.732 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.970 0.860 1.061 0.954 ;
      RECT 0.679 0.899 0.970 0.954 ;
      RECT 0.589 0.717 0.679 0.954 ;
      RECT 0.329 0.899 0.589 0.954 ;
      RECT 0.239 0.717 0.329 0.954 ;
  END
END AOI33X1

MACRO AOI32X4
  CLASS CORE ;
  FOREIGN AOI32X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.721 0.433 1.762 0.767 ;
      RECT 1.658 0.357 1.721 0.767 ;
      RECT 1.575 0.357 1.658 0.412 ;
      RECT 1.477 0.652 1.658 0.733 ;
      RECT 1.482 0.331 1.575 0.412 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.978 0.567 1.032 0.733 ;
      RECT 0.914 0.518 0.978 0.733 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.578 0.567 0.717 0.704 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.375 0.209 0.500 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.567 0.408 0.687 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.411 0.566 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.751 -0.080 1.800 0.080 ;
      RECT 1.658 -0.080 1.751 0.212 ;
      RECT 1.385 -0.080 1.658 0.080 ;
      RECT 1.323 -0.080 1.385 0.211 ;
      RECT 1.004 -0.080 1.323 0.080 ;
      RECT 0.911 -0.080 1.004 0.122 ;
      RECT 0.142 -0.080 0.911 0.080 ;
      RECT 0.049 -0.080 0.142 0.275 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.744 1.120 1.800 1.280 ;
      RECT 1.651 0.897 1.744 1.280 ;
      RECT 1.394 1.120 1.651 1.280 ;
      RECT 1.301 0.897 1.394 1.280 ;
      RECT 0.485 1.120 1.301 1.280 ;
      RECT 0.393 1.078 0.485 1.280 ;
      RECT 0.146 1.120 0.393 1.280 ;
      RECT 0.041 1.078 0.146 1.280 ;
      RECT 0.000 1.120 0.041 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.375 0.490 1.594 0.571 ;
      RECT 1.312 0.302 1.375 0.754 ;
      RECT 1.241 0.302 1.312 0.357 ;
      RECT 1.196 0.699 1.312 0.754 ;
      RECT 1.233 0.443 1.248 0.524 ;
      RECT 1.178 0.158 1.241 0.357 ;
      RECT 1.155 0.442 1.233 0.524 ;
      RECT 1.103 0.686 1.196 0.767 ;
      RECT 1.111 0.158 1.178 0.213 ;
      RECT 1.106 0.442 1.155 0.511 ;
      RECT 1.043 0.268 1.106 0.511 ;
      RECT 1.019 0.854 1.049 0.935 ;
      RECT 0.851 0.268 1.043 0.323 ;
      RECT 0.956 0.854 1.019 1.031 ;
      RECT 0.656 0.976 0.956 1.031 ;
      RECT 0.851 0.806 0.852 0.887 ;
      RECT 0.788 0.268 0.851 0.887 ;
      RECT 0.644 0.268 0.788 0.323 ;
      RECT 0.760 0.806 0.788 0.887 ;
      RECT 0.593 0.806 0.656 1.031 ;
      RECT 0.551 0.242 0.644 0.323 ;
      RECT 0.563 0.806 0.593 0.887 ;
      RECT 0.295 0.819 0.563 0.874 ;
      RECT 0.202 0.806 0.295 0.887 ;
  END
END AOI32X4

MACRO AOI32X1
  CLASS CORE ;
  FOREIGN AOI32X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.223 1.240 0.820 ;
      RECT 1.154 0.223 1.175 0.306 ;
      RECT 0.861 0.765 1.175 0.820 ;
      RECT 0.568 0.223 1.154 0.277 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.877 0.381 1.054 0.494 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.712 0.560 0.889 0.640 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.400 0.225 0.500 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.246 0.571 0.416 0.680 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.411 0.383 0.597 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 -0.080 1.300 0.080 ;
      RECT 0.948 -0.080 1.044 0.122 ;
      RECT 0.131 -0.080 0.948 0.080 ;
      RECT 0.066 -0.080 0.131 0.325 ;
      RECT 0.000 -0.080 0.066 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.552 1.120 1.300 1.280 ;
      RECT 0.456 0.925 0.552 1.280 ;
      RECT 0.146 1.120 0.456 1.280 ;
      RECT 0.051 0.800 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.739 0.908 1.159 0.963 ;
      RECT 0.674 0.800 0.739 0.963 ;
      RECT 0.253 0.800 0.674 0.855 ;
  END
END AOI32X1

MACRO AOI31XL
  CLASS CORE ;
  FOREIGN AOI31XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.836 0.280 0.841 0.361 ;
      RECT 0.773 0.280 0.836 0.790 ;
      RECT 0.551 0.280 0.773 0.335 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.642 0.565 0.705 0.656 ;
      RECT 0.535 0.567 0.642 0.656 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.381 0.142 0.520 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.567 0.405 0.650 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.420 0.390 0.622 0.500 ;
      RECT 0.419 0.439 0.420 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.836 -0.080 0.900 0.080 ;
      RECT 0.743 -0.080 0.836 0.122 ;
      RECT 0.142 -0.080 0.743 0.080 ;
      RECT 0.049 -0.080 0.142 0.275 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.502 1.120 0.900 1.280 ;
      RECT 0.409 1.078 0.502 1.280 ;
      RECT 0.149 1.120 0.409 1.280 ;
      RECT 0.048 1.078 0.149 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.202 0.760 0.655 0.840 ;
  END
END AOI31XL

MACRO AOI31X1
  CLASS CORE ;
  FOREIGN AOI31X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.825 0.201 0.841 0.756 ;
      RECT 0.779 0.201 0.825 0.958 ;
      RECT 0.758 0.201 0.779 0.367 ;
      RECT 0.762 0.701 0.779 0.958 ;
      RECT 0.551 0.201 0.758 0.256 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.715 0.501 0.716 0.583 ;
      RECT 0.608 0.501 0.715 0.633 ;
      RECT 0.578 0.567 0.608 0.633 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.420 0.142 0.571 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.218 0.558 0.353 0.668 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.398 0.529 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.122 ;
      RECT 0.142 -0.080 0.758 0.080 ;
      RECT 0.049 -0.080 0.142 0.198 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.491 1.120 0.900 1.280 ;
      RECT 0.398 0.915 0.491 1.280 ;
      RECT 0.142 1.120 0.398 1.280 ;
      RECT 0.049 0.916 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.224 0.724 0.665 0.779 ;
  END
END AOI31X1

MACRO AOI2BB2X4
  CLASS CORE ;
  FOREIGN AOI2BB2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.117 0.167 2.217 0.500 ;
      RECT 0.928 0.269 2.117 0.324 ;
      RECT 0.924 0.979 1.245 1.033 ;
      RECT 0.924 0.221 0.928 0.324 ;
      RECT 0.864 0.221 0.924 1.033 ;
      RECT 0.819 0.979 0.864 1.033 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.013 0.587 2.295 0.642 ;
      RECT 1.953 0.438 2.013 0.642 ;
      RECT 1.330 0.438 1.953 0.493 ;
      RECT 1.181 0.438 1.330 0.494 ;
      RECT 1.120 0.438 1.181 0.554 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.564 0.567 1.697 0.668 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.563 0.706 0.637 0.761 ;
      RECT 0.503 0.460 0.563 0.992 ;
      RECT 0.137 0.937 0.503 0.992 ;
      RECT 0.125 0.894 0.137 0.992 ;
      RECT 0.064 0.562 0.125 0.992 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.197 0.408 0.320 0.526 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.863 -0.080 2.600 0.080 ;
      RECT 1.774 -0.080 1.863 0.198 ;
      RECT 1.132 -0.080 1.774 0.080 ;
      RECT 1.043 -0.080 1.132 0.198 ;
      RECT 0.653 -0.080 1.043 0.080 ;
      RECT 0.563 -0.080 0.653 0.122 ;
      RECT 0.240 -0.080 0.563 0.080 ;
      RECT 0.151 -0.080 0.240 0.198 ;
      RECT 0.000 -0.080 0.151 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.253 1.120 2.600 1.280 ;
      RECT 2.164 0.980 2.253 1.280 ;
      RECT 1.917 1.120 2.164 1.280 ;
      RECT 1.828 0.980 1.917 1.280 ;
      RECT 1.581 1.120 1.828 1.280 ;
      RECT 1.492 0.980 1.581 1.280 ;
      RECT 0.725 1.120 1.492 1.280 ;
      RECT 0.636 1.078 0.725 1.280 ;
      RECT 0.137 1.120 0.636 1.280 ;
      RECT 0.047 1.078 0.137 1.280 ;
      RECT 0.000 1.120 0.047 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.987 0.737 2.421 0.792 ;
      RECT 0.742 0.270 0.802 0.538 ;
      RECT 0.441 0.270 0.742 0.325 ;
      RECT 0.381 0.270 0.441 0.785 ;
      RECT 0.358 0.270 0.381 0.325 ;
      RECT 0.356 0.698 0.381 0.785 ;
  END
END AOI2BB2X4

MACRO AOI2BB2X2
  CLASS CORE ;
  FOREIGN AOI2BB2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.508 0.306 1.542 0.361 ;
      RECT 1.446 0.192 1.508 0.977 ;
      RECT 0.773 0.192 1.446 0.246 ;
      RECT 1.304 0.923 1.446 0.977 ;
      RECT 1.203 0.923 1.304 1.040 ;
      RECT 1.187 0.967 1.203 1.040 ;
      RECT 1.094 0.986 1.187 1.040 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.104 0.543 1.201 0.737 ;
      RECT 0.512 0.682 1.104 0.737 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.294 0.379 1.371 0.498 ;
      RECT 0.672 0.379 1.294 0.433 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.343 0.388 0.496 0.500 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.445 0.140 0.633 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.072 -0.080 1.600 0.080 ;
      RECT 0.980 -0.080 1.072 0.122 ;
      RECT 0.516 -0.080 0.980 0.080 ;
      RECT 0.424 -0.080 0.516 0.289 ;
      RECT 0.140 -0.080 0.424 0.080 ;
      RECT 0.048 -0.080 0.140 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 1.120 1.600 1.280 ;
      RECT 1.449 1.078 1.541 1.280 ;
      RECT 0.840 1.120 1.449 1.280 ;
      RECT 0.749 0.988 0.840 1.280 ;
      RECT 0.496 1.120 0.749 1.280 ;
      RECT 0.404 0.988 0.496 1.280 ;
      RECT 0.000 1.120 0.404 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.576 0.808 1.358 0.863 ;
      RECT 0.276 0.571 0.991 0.626 ;
      RECT 0.214 0.288 0.276 0.788 ;
      RECT 0.048 0.733 0.214 0.788 ;
  END
END AOI2BB2X2

MACRO AOI2BB2X1
  CLASS CORE ;
  FOREIGN AOI2BB2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.097 0.265 1.162 1.049 ;
      RECT 0.760 0.265 1.097 0.320 ;
      RECT 0.989 0.567 1.097 0.633 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.550 0.661 0.703 0.767 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.803 0.536 0.868 0.627 ;
      RECT 0.737 0.536 0.803 0.590 ;
      RECT 0.673 0.501 0.737 0.590 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.053 0.433 0.134 0.620 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.224 0.536 0.348 0.651 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.069 -0.080 1.300 0.080 ;
      RECT 0.974 -0.080 1.069 0.122 ;
      RECT 0.484 -0.080 0.974 0.080 ;
      RECT 0.388 -0.080 0.484 0.122 ;
      RECT 0.146 -0.080 0.388 0.080 ;
      RECT 0.051 -0.080 0.146 0.122 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.816 1.120 1.300 1.280 ;
      RECT 0.720 0.989 0.816 1.280 ;
      RECT 0.146 1.120 0.720 1.280 ;
      RECT 0.051 1.078 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.644 0.821 0.996 0.876 ;
      RECT 0.910 0.375 0.975 0.474 ;
      RECT 0.478 0.375 0.910 0.430 ;
      RECT 0.580 0.821 0.644 1.042 ;
      RECT 0.518 0.987 0.580 1.042 ;
      RECT 0.414 0.375 0.478 0.814 ;
      RECT 0.300 0.375 0.414 0.430 ;
      RECT 0.381 0.726 0.414 0.814 ;
      RECT 0.235 0.313 0.300 0.430 ;
  END
END AOI2BB2X1

MACRO AOI2BB1XL
  CLASS CORE ;
  FOREIGN AOI2BB1XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.792 0.839 0.841 0.894 ;
      RECT 0.730 0.386 0.792 0.907 ;
      RECT 0.574 0.386 0.730 0.440 ;
      RECT 0.511 0.348 0.574 0.440 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.636 0.532 0.767 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.147 0.538 0.301 0.627 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.048 0.689 0.199 0.789 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.346 -0.080 0.900 0.080 ;
      RECT 0.254 -0.080 0.346 0.122 ;
      RECT 0.000 -0.080 0.254 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.447 1.120 0.900 1.280 ;
      RECT 0.355 1.078 0.447 1.280 ;
      RECT 0.000 1.120 0.355 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.595 0.496 0.657 0.901 ;
      RECT 0.447 0.496 0.595 0.551 ;
      RECT 0.049 0.846 0.595 0.901 ;
      RECT 0.385 0.313 0.447 0.551 ;
      RECT 0.123 0.313 0.385 0.368 ;
  END
END AOI2BB1XL

MACRO AOI2BB1X1
  CLASS CORE ;
  FOREIGN AOI2BB1X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.794 0.292 0.841 0.761 ;
      RECT 0.779 0.292 0.794 0.986 ;
      RECT 0.570 0.292 0.779 0.346 ;
      RECT 0.731 0.706 0.779 0.986 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.535 0.665 0.536 0.761 ;
      RECT 0.359 0.665 0.535 0.767 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.150 0.424 0.322 0.505 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.567 0.218 0.679 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.346 -0.080 0.900 0.080 ;
      RECT 0.254 -0.080 0.346 0.122 ;
      RECT 0.000 -0.080 0.254 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.447 1.120 0.900 1.280 ;
      RECT 0.355 1.078 0.447 1.280 ;
      RECT 0.000 1.120 0.355 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.663 0.501 0.715 0.587 ;
      RECT 0.600 0.446 0.663 0.894 ;
      RECT 0.462 0.446 0.600 0.501 ;
      RECT 0.049 0.839 0.600 0.894 ;
      RECT 0.400 0.311 0.462 0.501 ;
      RECT 0.123 0.311 0.400 0.365 ;
  END
END AOI2BB1X1

MACRO AOI22XL
  CLASS CORE ;
  FOREIGN AOI22XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.282 0.862 0.815 ;
      RECT 0.779 0.282 0.799 0.361 ;
      RECT 0.665 0.761 0.799 0.815 ;
      RECT 0.502 0.282 0.779 0.337 ;
      RECT 0.573 0.748 0.665 0.829 ;
      RECT 0.409 0.269 0.502 0.350 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.396 0.169 0.511 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.325 0.560 0.417 0.649 ;
      RECT 0.218 0.567 0.325 0.649 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.716 0.571 0.731 0.652 ;
      RECT 0.567 0.562 0.716 0.652 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.601 0.425 0.603 0.500 ;
      RECT 0.481 0.412 0.601 0.500 ;
      RECT 0.417 0.425 0.481 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.840 -0.080 0.900 0.080 ;
      RECT 0.747 -0.080 0.840 0.122 ;
      RECT 0.142 -0.080 0.747 0.080 ;
      RECT 0.049 -0.080 0.142 0.122 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.176 1.120 0.900 1.280 ;
      RECT 0.063 1.078 0.176 1.280 ;
      RECT 0.000 1.120 0.063 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.453 0.994 0.821 1.049 ;
      RECT 0.390 0.762 0.453 1.049 ;
      RECT 0.142 0.762 0.390 0.817 ;
      RECT 0.049 0.749 0.142 0.830 ;
  END
END AOI22XL

MACRO AOI22X4
  CLASS CORE ;
  FOREIGN AOI22X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.284 0.439 2.346 0.985 ;
      RECT 2.263 0.300 2.284 0.633 ;
      RECT 2.024 0.930 2.284 0.985 ;
      RECT 2.181 0.287 2.263 0.633 ;
      RECT 0.049 0.287 2.181 0.342 ;
      RECT 1.939 0.930 2.024 1.033 ;
      RECT 1.905 0.967 1.939 1.033 ;
      RECT 1.261 0.979 1.905 1.033 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.066 0.438 1.081 0.493 ;
      RECT 1.004 0.438 1.066 0.494 ;
      RECT 0.237 0.439 1.004 0.494 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.656 0.587 0.770 0.642 ;
      RECT 0.594 0.573 0.656 0.642 ;
      RECT 0.114 0.587 0.594 0.642 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.288 0.439 1.872 0.494 ;
      RECT 1.247 0.439 1.288 0.500 ;
      RECT 1.185 0.439 1.247 0.654 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.043 0.504 2.105 0.627 ;
      RECT 1.370 0.573 2.043 0.627 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.872 -0.080 2.500 0.080 ;
      RECT 1.780 -0.080 1.872 0.203 ;
      RECT 1.180 -0.080 1.780 0.080 ;
      RECT 1.088 -0.080 1.180 0.203 ;
      RECT 0.487 -0.080 1.088 0.080 ;
      RECT 0.395 -0.080 0.487 0.203 ;
      RECT 0.000 -0.080 0.395 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.006 1.120 2.500 1.280 ;
      RECT 0.915 0.980 1.006 1.280 ;
      RECT 0.660 1.120 0.915 1.280 ;
      RECT 0.568 0.980 0.660 1.280 ;
      RECT 0.314 1.120 0.568 1.280 ;
      RECT 0.222 0.980 0.314 1.280 ;
      RECT 0.000 1.120 0.222 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.049 0.737 2.219 0.792 ;
  END
END AOI22X4

MACRO AOI22X2
  CLASS CORE ;
  FOREIGN AOI22X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.321 1.542 0.761 ;
      RECT 0.393 0.321 1.480 0.376 ;
      RECT 1.368 0.706 1.480 0.761 ;
      RECT 1.302 0.706 1.368 0.789 ;
      RECT 0.932 0.735 1.302 0.789 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.653 0.456 0.715 0.575 ;
      RECT 0.298 0.456 0.653 0.511 ;
      RECT 0.246 0.439 0.298 0.511 ;
      RECT 0.185 0.439 0.246 0.562 ;
      RECT 0.113 0.493 0.185 0.562 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.329 0.573 0.475 0.663 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.356 0.438 1.418 0.551 ;
      RECT 1.009 0.438 1.356 0.493 ;
      RECT 0.944 0.438 1.009 0.494 ;
      RECT 0.882 0.438 0.944 0.664 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.061 0.567 1.207 0.661 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.444 -0.080 1.600 0.080 ;
      RECT 1.352 -0.080 1.444 0.122 ;
      RECT 0.787 -0.080 1.352 0.080 ;
      RECT 0.695 -0.080 0.787 0.122 ;
      RECT 0.140 -0.080 0.695 0.080 ;
      RECT 0.048 -0.080 0.140 0.305 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.657 1.120 1.600 1.280 ;
      RECT 0.566 0.888 0.657 1.280 ;
      RECT 0.312 1.120 0.566 1.280 ;
      RECT 0.221 0.888 0.312 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.815 0.886 1.541 0.940 ;
      RECT 0.815 0.732 0.830 0.787 ;
      RECT 0.753 0.732 0.815 0.940 ;
      RECT 0.048 0.732 0.753 0.787 ;
  END
END AOI22X2

MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.265 0.862 0.754 ;
      RECT 0.779 0.265 0.799 0.361 ;
      RECT 0.676 0.699 0.799 0.754 ;
      RECT 0.491 0.265 0.779 0.320 ;
      RECT 0.584 0.699 0.676 0.780 ;
      RECT 0.398 0.252 0.491 0.333 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.052 0.421 0.145 0.589 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.239 0.567 0.415 0.663 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.577 0.538 0.731 0.633 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.499 0.394 0.592 0.475 ;
      RECT 0.481 0.407 0.499 0.475 ;
      RECT 0.419 0.407 0.481 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.122 ;
      RECT 0.142 -0.080 0.758 0.080 ;
      RECT 0.049 -0.080 0.142 0.330 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.322 1.120 0.900 1.280 ;
      RECT 0.229 1.078 0.322 1.280 ;
      RECT 0.000 1.120 0.229 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.758 0.854 0.851 0.935 ;
      RECT 0.502 0.880 0.758 0.935 ;
      RECT 0.409 0.865 0.502 0.946 ;
      RECT 0.142 0.879 0.409 0.933 ;
      RECT 0.049 0.726 0.142 0.933 ;
  END
END AOI22X1

MACRO AOI222XL
  CLASS CORE ;
  FOREIGN AOI222XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.282 0.270 1.343 0.737 ;
      RECT 0.048 0.270 1.282 0.325 ;
      RECT 1.262 0.627 1.282 0.737 ;
      RECT 1.051 0.682 1.262 0.737 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.568 0.337 0.687 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.433 0.138 0.564 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.404 0.411 0.550 0.500 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.688 0.433 0.834 0.524 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.106 0.439 1.198 0.605 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.921 0.392 1.022 0.523 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.286 -0.080 1.400 0.080 ;
      RECT 1.196 -0.080 1.286 0.122 ;
      RECT 0.500 -0.080 1.196 0.080 ;
      RECT 0.410 -0.080 0.500 0.200 ;
      RECT 0.000 -0.080 0.410 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.308 1.120 1.400 1.280 ;
      RECT 0.217 1.065 0.308 1.280 ;
      RECT 0.000 1.120 0.217 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.552 0.987 1.290 1.042 ;
      RECT 0.196 0.801 0.790 0.856 ;
  END
END AOI222XL

MACRO AOI222X1
  CLASS CORE ;
  FOREIGN AOI222X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.282 0.281 1.343 0.743 ;
      RECT 0.048 0.281 1.282 0.336 ;
      RECT 1.083 0.688 1.282 0.743 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.232 0.405 0.380 0.507 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.439 0.122 0.633 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.506 0.586 0.627 ;
      RECT 0.407 0.573 0.488 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.701 0.433 0.838 0.535 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.087 0.433 1.188 0.587 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.912 0.444 1.013 0.627 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.269 -0.080 1.400 0.080 ;
      RECT 1.179 -0.080 1.269 0.122 ;
      RECT 0.508 -0.080 1.179 0.080 ;
      RECT 0.418 -0.080 0.508 0.122 ;
      RECT 0.000 -0.080 0.418 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.477 1.120 1.400 1.280 ;
      RECT 0.387 0.917 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.941 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.574 0.910 1.343 0.964 ;
      RECT 0.707 0.685 0.834 0.739 ;
      RECT 0.646 0.685 0.707 0.817 ;
      RECT 0.217 0.762 0.646 0.817 ;
  END
END AOI222X1

MACRO AOI221XL
  CLASS CORE ;
  FOREIGN AOI221XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.236 1.240 0.743 ;
      RECT 1.154 0.236 1.175 0.306 ;
      RECT 1.092 0.688 1.175 0.743 ;
      RECT 0.612 0.236 1.154 0.290 ;
      RECT 0.547 0.161 0.612 0.290 ;
      RECT 0.497 0.161 0.547 0.233 ;
      RECT 0.411 0.161 0.497 0.215 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.019 0.573 1.054 0.627 ;
      RECT 0.954 0.433 1.019 0.627 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.313 0.146 0.500 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.225 0.562 0.377 0.671 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.722 0.374 0.868 0.494 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.439 0.553 0.613 ;
      RECT 0.432 0.439 0.488 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.878 -0.080 1.300 0.080 ;
      RECT 0.782 -0.080 0.878 0.122 ;
      RECT 0.146 -0.080 0.782 0.080 ;
      RECT 0.051 -0.080 0.146 0.198 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.461 1.120 1.300 1.280 ;
      RECT 0.366 1.078 0.461 1.280 ;
      RECT 0.146 1.120 0.366 1.280 ;
      RECT 0.051 1.078 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.563 0.995 0.974 1.050 ;
      RECT 0.720 0.671 0.816 0.867 ;
      RECT 0.304 0.812 0.720 0.867 ;
      RECT 0.208 0.740 0.304 0.936 ;
  END
END AOI221XL

MACRO AOI221X2
  CLASS CORE ;
  FOREIGN AOI221X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.807 0.312 1.868 0.836 ;
      RECT 1.457 0.312 1.807 0.367 ;
      RECT 1.761 0.755 1.807 0.836 ;
      RECT 1.391 0.300 1.457 0.367 ;
      RECT 1.330 0.225 1.391 0.367 ;
      RECT 0.387 0.225 1.330 0.280 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.678 0.439 1.739 0.543 ;
      RECT 1.457 0.439 1.678 0.494 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.663 0.493 0.711 0.558 ;
      RECT 0.562 0.433 0.663 0.558 ;
      RECT 0.077 0.504 0.562 0.558 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 0.375 0.414 0.430 ;
      RECT 0.212 0.306 0.313 0.430 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.993 0.595 1.572 0.650 ;
      RECT 0.932 0.573 0.993 0.650 ;
      RECT 0.917 0.595 0.932 0.650 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.087 0.396 1.233 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.636 -0.080 2.100 0.080 ;
      RECT 1.546 -0.080 1.636 0.198 ;
      RECT 0.870 -0.080 1.546 0.080 ;
      RECT 0.780 -0.080 0.870 0.122 ;
      RECT 0.138 -0.080 0.780 0.080 ;
      RECT 0.048 -0.080 0.138 0.198 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.817 1.120 2.100 1.280 ;
      RECT 0.727 0.903 0.817 1.280 ;
      RECT 0.477 1.120 0.727 1.280 ;
      RECT 0.387 0.903 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.903 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.912 0.962 2.020 1.017 ;
      RECT 0.944 0.768 1.511 0.823 ;
      RECT 0.883 0.707 0.944 0.823 ;
      RECT 0.217 0.707 0.883 0.762 ;
  END
END AOI221X2

MACRO AOI221X1
  CLASS CORE ;
  FOREIGN AOI221X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.257 1.240 0.761 ;
      RECT 0.703 0.257 1.175 0.312 ;
      RECT 1.165 0.627 1.175 0.754 ;
      RECT 0.696 0.227 0.703 0.312 ;
      RECT 0.632 0.189 0.696 0.312 ;
      RECT 0.411 0.189 0.632 0.244 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 0.573 1.054 0.627 ;
      RECT 0.979 0.393 1.044 0.627 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.049 0.306 0.146 0.461 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.225 0.520 0.380 0.633 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.803 0.379 0.868 0.494 ;
      RECT 0.667 0.379 0.803 0.433 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.432 0.306 0.560 0.431 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.878 -0.080 1.300 0.080 ;
      RECT 0.782 -0.080 0.878 0.122 ;
      RECT 0.146 -0.080 0.782 0.080 ;
      RECT 0.051 -0.080 0.146 0.229 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.506 1.120 1.300 1.280 ;
      RECT 0.411 0.916 0.506 1.280 ;
      RECT 0.146 1.120 0.411 1.280 ;
      RECT 0.051 0.916 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.609 0.862 1.065 0.917 ;
      RECT 0.231 0.689 0.885 0.744 ;
  END
END AOI221X1

MACRO AOI21XL
  CLASS CORE ;
  FOREIGN AOI21XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.634 0.295 0.643 0.627 ;
      RECT 0.582 0.295 0.634 0.830 ;
      RECT 0.387 0.295 0.582 0.350 ;
      RECT 0.573 0.573 0.582 0.830 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.362 0.411 0.513 0.500 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.045 0.417 0.138 0.562 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.567 0.379 0.662 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.626 -0.080 0.700 0.080 ;
      RECT 0.536 -0.080 0.626 0.122 ;
      RECT 0.138 -0.080 0.536 0.080 ;
      RECT 0.048 -0.080 0.138 0.331 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.223 1.078 0.313 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.435 0.995 0.498 1.050 ;
      RECT 0.374 0.952 0.435 1.050 ;
      RECT 0.123 0.952 0.374 1.007 ;
      RECT 0.062 0.749 0.123 1.007 ;
  END
END AOI21XL

MACRO AOI21X4
  CLASS CORE ;
  FOREIGN AOI21X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.668 0.896 1.713 0.977 ;
      RECT 1.620 0.579 1.668 0.977 ;
      RECT 1.605 0.579 1.620 0.964 ;
      RECT 1.582 0.579 1.605 0.633 ;
      RECT 1.364 0.910 1.605 0.964 ;
      RECT 1.478 0.300 1.582 0.633 ;
      RECT 1.319 0.337 1.478 0.392 ;
      RECT 1.271 0.896 1.364 0.977 ;
      RECT 1.208 0.274 1.319 0.392 ;
      RECT 0.049 0.274 1.208 0.329 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.238 0.496 1.402 0.635 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.068 0.452 1.098 0.533 ;
      RECT 1.005 0.392 1.068 0.533 ;
      RECT 0.661 0.392 1.005 0.446 ;
      RECT 0.492 0.392 0.661 0.494 ;
      RECT 0.415 0.392 0.492 0.507 ;
      RECT 0.400 0.426 0.415 0.507 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.807 0.573 0.841 0.627 ;
      RECT 0.745 0.530 0.807 0.627 ;
      RECT 0.218 0.570 0.745 0.625 ;
      RECT 0.207 0.567 0.218 0.625 ;
      RECT 0.145 0.469 0.207 0.625 ;
      RECT 0.115 0.469 0.145 0.574 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.550 -0.080 1.800 0.080 ;
      RECT 1.458 -0.080 1.550 0.122 ;
      RECT 1.190 -0.080 1.458 0.080 ;
      RECT 1.098 -0.080 1.190 0.198 ;
      RECT 0.492 -0.080 1.098 0.080 ;
      RECT 0.400 -0.080 0.492 0.198 ;
      RECT 0.000 -0.080 0.400 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.015 1.120 1.800 1.280 ;
      RECT 0.922 0.941 1.015 1.280 ;
      RECT 0.665 1.120 0.922 1.280 ;
      RECT 0.573 0.941 0.665 1.280 ;
      RECT 0.316 1.120 0.573 1.280 ;
      RECT 0.224 0.941 0.316 1.280 ;
      RECT 0.000 1.120 0.224 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.049 0.698 1.538 0.752 ;
  END
END AOI21X4

MACRO AOI21X2
  CLASS CORE ;
  FOREIGN AOI21X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.030 0.345 1.095 0.789 ;
      RECT 0.867 0.345 1.030 0.400 ;
      RECT 0.989 0.706 1.030 0.789 ;
      RECT 0.974 0.735 0.989 0.789 ;
      RECT 0.771 0.268 0.867 0.400 ;
      RECT 0.300 0.345 0.771 0.400 ;
      RECT 0.235 0.294 0.300 0.400 ;
      RECT 0.146 0.294 0.235 0.349 ;
      RECT 0.051 0.268 0.146 0.349 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.830 0.485 0.936 0.627 ;
      RECT 0.803 0.573 0.830 0.627 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.311 0.595 0.518 0.669 ;
      RECT 0.246 0.573 0.311 0.669 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.146 0.457 0.763 0.512 ;
      RECT 0.039 0.433 0.146 0.530 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.082 -0.080 1.300 0.080 ;
      RECT 0.986 -0.080 1.082 0.122 ;
      RECT 0.506 -0.080 0.986 0.080 ;
      RECT 0.411 -0.080 0.506 0.275 ;
      RECT 0.000 -0.080 0.411 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.687 1.120 1.300 1.280 ;
      RECT 0.591 0.888 0.687 1.280 ;
      RECT 0.326 1.120 0.591 1.280 ;
      RECT 0.231 0.888 0.326 1.280 ;
      RECT 0.000 1.120 0.231 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.154 0.873 1.249 0.954 ;
      RECT 0.871 0.873 1.154 0.927 ;
      RECT 0.806 0.732 0.871 0.927 ;
      RECT 0.051 0.732 0.806 0.787 ;
  END
END AOI21X2

MACRO AOI21X1
  CLASS CORE ;
  FOREIGN AOI21X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.603 0.321 0.664 0.940 ;
      RECT 0.477 0.321 0.603 0.376 ;
      RECT 0.582 0.706 0.603 0.940 ;
      RECT 0.557 0.860 0.582 0.940 ;
      RECT 0.387 0.295 0.477 0.376 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.477 0.439 0.542 0.627 ;
      RECT 0.407 0.439 0.477 0.494 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.138 0.492 0.141 0.615 ;
      RECT 0.050 0.433 0.138 0.615 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.293 0.568 0.379 0.623 ;
      RECT 0.232 0.306 0.293 0.623 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.626 -0.080 0.700 0.080 ;
      RECT 0.536 -0.080 0.626 0.122 ;
      RECT 0.138 -0.080 0.536 0.080 ;
      RECT 0.048 -0.080 0.138 0.334 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.308 1.120 0.700 1.280 ;
      RECT 0.217 0.852 0.308 1.280 ;
      RECT 0.000 1.120 0.217 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.048 0.696 0.477 0.751 ;
  END
END AOI21X1

MACRO AND4X4
  CLASS CORE ;
  FOREIGN AND4X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.759 0.567 1.780 0.900 ;
      RECT 1.696 0.356 1.759 0.900 ;
      RECT 1.676 0.331 1.696 0.900 ;
      RECT 1.675 0.331 1.676 0.439 ;
      RECT 1.675 0.567 1.676 0.900 ;
      RECT 1.570 0.331 1.675 0.412 ;
      RECT 1.532 0.815 1.675 0.900 ;
      RECT 1.438 0.815 1.532 1.039 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.328 0.439 1.364 0.494 ;
      RECT 1.264 0.439 1.328 0.650 ;
      RECT 1.213 0.567 1.264 0.650 ;
      RECT 1.178 0.595 1.213 0.650 ;
      RECT 1.114 0.595 1.178 0.888 ;
      RECT 0.145 0.833 1.114 0.888 ;
      RECT 0.145 0.640 0.146 0.767 ;
      RECT 0.081 0.640 0.145 0.888 ;
      RECT 0.039 0.640 0.081 0.767 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.988 0.379 1.051 0.721 ;
      RECT 0.948 0.379 0.988 0.439 ;
      RECT 0.344 0.379 0.948 0.433 ;
      RECT 0.344 0.539 0.364 0.636 ;
      RECT 0.281 0.379 0.344 0.636 ;
      RECT 0.220 0.493 0.281 0.636 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.766 0.489 0.871 0.629 ;
      RECT 0.460 0.489 0.766 0.544 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.579 0.625 0.689 0.773 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.862 -0.080 2.000 0.080 ;
      RECT 1.769 -0.080 1.862 0.211 ;
      RECT 1.466 -0.080 1.769 0.080 ;
      RECT 1.372 -0.080 1.466 0.250 ;
      RECT 0.143 -0.080 1.372 0.080 ;
      RECT 0.050 -0.080 0.143 0.334 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.751 1.120 2.000 1.280 ;
      RECT 1.643 1.078 1.751 1.280 ;
      RECT 1.225 1.120 1.643 1.280 ;
      RECT 1.131 1.078 1.225 1.280 ;
      RECT 0.782 1.120 1.131 1.280 ;
      RECT 0.689 1.078 0.782 1.280 ;
      RECT 0.358 1.120 0.689 1.280 ;
      RECT 0.251 1.078 0.358 1.280 ;
      RECT 0.000 1.120 0.251 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.507 0.507 1.574 0.588 ;
      RECT 1.444 0.329 1.507 0.761 ;
      RECT 1.227 0.329 1.444 0.383 ;
      RECT 1.306 0.706 1.444 0.761 ;
      RECT 1.242 0.706 1.306 0.999 ;
      RECT 0.999 0.944 1.242 0.999 ;
      RECT 1.164 0.254 1.227 0.383 ;
      RECT 0.804 0.254 1.164 0.308 ;
      RECT 0.905 0.944 0.999 1.039 ;
      RECT 0.573 0.944 0.905 0.999 ;
      RECT 0.711 0.240 0.804 0.321 ;
      RECT 0.479 0.944 0.573 1.039 ;
  END
END AND4X4

MACRO AND4X2
  CLASS CORE ;
  FOREIGN AND4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.049 0.700 1.061 0.767 ;
      RECT 1.031 0.358 1.049 0.767 ;
      RECT 0.985 0.199 1.031 0.964 ;
      RECT 0.967 0.199 0.985 0.413 ;
      RECT 0.967 0.648 0.985 0.964 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.694 0.524 0.733 0.606 ;
      RECT 0.610 0.439 0.694 0.606 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.478 0.581 0.542 0.761 ;
      RECT 0.426 0.706 0.478 0.761 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.279 0.537 0.358 0.646 ;
      RECT 0.222 0.537 0.279 0.645 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.398 0.157 0.556 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.815 -0.080 1.100 0.080 ;
      RECT 0.721 -0.080 0.815 0.122 ;
      RECT 0.000 -0.080 0.721 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.838 1.120 1.100 1.280 ;
      RECT 0.724 1.064 0.838 1.280 ;
      RECT 0.514 1.120 0.724 1.280 ;
      RECT 0.419 1.078 0.514 1.280 ;
      RECT 0.158 1.120 0.419 1.280 ;
      RECT 0.049 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.889 0.473 0.919 0.556 ;
      RECT 0.825 0.211 0.889 0.889 ;
      RECT 0.156 0.211 0.825 0.265 ;
      RECT 0.208 0.835 0.825 0.889 ;
      RECT 0.076 0.211 0.156 0.343 ;
      RECT 0.061 0.250 0.076 0.343 ;
  END
END AND4X2

MACRO AND4X1
  CLASS CORE ;
  FOREIGN AND4X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.044 0.761 1.061 0.905 ;
      RECT 0.981 0.244 1.044 0.905 ;
      RECT 0.950 0.244 0.981 0.325 ;
      RECT 0.956 0.761 0.981 0.905 ;
      RECT 0.950 0.800 0.956 0.905 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.703 0.573 0.857 0.696 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.392 0.567 0.511 0.696 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.175 0.399 0.328 0.545 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.615 0.147 0.776 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.833 -0.080 1.100 0.080 ;
      RECT 0.739 -0.080 0.833 0.122 ;
      RECT 0.000 -0.080 0.739 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.861 1.120 1.100 1.280 ;
      RECT 0.258 1.078 0.861 1.280 ;
      RECT 0.000 1.120 0.258 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.878 0.401 0.908 0.482 ;
      RECT 0.814 0.223 0.878 0.482 ;
      RECT 0.144 0.223 0.814 0.277 ;
      RECT 0.639 0.414 0.814 0.469 ;
      RECT 0.628 0.414 0.639 0.824 ;
      RECT 0.575 0.414 0.628 0.887 ;
      RECT 0.533 0.751 0.575 0.887 ;
      RECT 0.144 0.832 0.533 0.887 ;
      RECT 0.050 0.223 0.144 0.304 ;
  END
END AND4X1

MACRO AOI211XL
  CLASS CORE ;
  FOREIGN AOI211XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.799 0.274 0.862 0.761 ;
      RECT 0.398 0.274 0.799 0.329 ;
      RECT 0.758 0.706 0.799 0.761 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.412 0.555 0.580 0.645 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.674 0.433 0.736 0.592 ;
      RECT 0.577 0.433 0.674 0.500 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.465 0.142 0.633 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.217 0.393 0.375 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.671 -0.080 0.900 0.080 ;
      RECT 0.578 -0.080 0.671 0.122 ;
      RECT 0.142 -0.080 0.578 0.080 ;
      RECT 0.049 -0.080 0.142 0.280 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.295 1.120 0.900 1.280 ;
      RECT 0.202 1.078 0.295 1.280 ;
      RECT 0.000 1.120 0.202 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.049 0.704 0.502 0.758 ;
  END
END AOI211XL

MACRO AOI211X2
  CLASS CORE ;
  FOREIGN AOI211X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.471 0.249 1.533 0.761 ;
      RECT 1.414 0.249 1.471 0.304 ;
      RECT 1.177 0.706 1.471 0.761 ;
      RECT 1.323 0.223 1.414 0.304 ;
      RECT 0.980 0.236 1.323 0.290 ;
      RECT 1.100 0.706 1.177 0.807 ;
      RECT 1.086 0.726 1.100 0.807 ;
      RECT 0.762 0.223 0.980 0.304 ;
      RECT 0.749 0.223 0.762 0.290 ;
      RECT 0.143 0.236 0.749 0.290 ;
      RECT 0.051 0.223 0.143 0.304 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.345 0.365 1.407 0.539 ;
      RECT 1.282 0.365 1.345 0.439 ;
      RECT 0.905 0.365 1.282 0.420 ;
      RECT 0.843 0.365 0.905 0.627 ;
      RECT 0.769 0.550 0.843 0.627 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.021 0.550 1.207 0.645 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.236 0.539 0.399 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.601 0.494 0.615 0.621 ;
      RECT 0.539 0.399 0.601 0.621 ;
      RECT 0.207 0.399 0.539 0.454 ;
      RECT 0.524 0.540 0.539 0.621 ;
      RECT 0.120 0.386 0.207 0.467 ;
      RECT 0.116 0.386 0.120 0.494 ;
      RECT 0.058 0.399 0.116 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.208 -0.080 1.600 0.080 ;
      RECT 1.116 -0.080 1.208 0.122 ;
      RECT 0.498 -0.080 1.116 0.080 ;
      RECT 0.407 -0.080 0.498 0.122 ;
      RECT 0.000 -0.080 0.407 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.659 1.120 1.600 1.280 ;
      RECT 0.567 0.925 0.659 1.280 ;
      RECT 0.314 1.120 0.567 1.280 ;
      RECT 0.222 0.925 0.314 1.280 ;
      RECT 0.000 1.120 0.222 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.430 0.881 1.522 0.962 ;
      RECT 0.937 0.894 1.430 0.949 ;
      RECT 0.875 0.688 0.937 0.949 ;
      RECT 0.050 0.688 0.875 0.743 ;
  END
END AOI211X2

MACRO AOI211X1
  CLASS CORE ;
  FOREIGN AOI211X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.840 0.261 0.867 0.761 ;
      RECT 0.821 0.261 0.840 0.975 ;
      RECT 0.805 0.192 0.821 0.975 ;
      RECT 0.758 0.192 0.805 0.342 ;
      RECT 0.747 0.661 0.805 0.975 ;
      RECT 0.500 0.192 0.758 0.246 ;
      RECT 0.438 0.192 0.500 0.329 ;
      RECT 0.398 0.274 0.438 0.329 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.515 0.558 0.633 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.685 0.436 0.742 0.536 ;
      RECT 0.679 0.436 0.685 0.761 ;
      RECT 0.622 0.481 0.679 0.761 ;
      RECT 0.599 0.706 0.622 0.761 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.524 0.176 0.645 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.322 0.400 0.390 0.455 ;
      RECT 0.239 0.306 0.322 0.455 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.640 -0.080 0.900 0.080 ;
      RECT 0.547 -0.080 0.640 0.122 ;
      RECT 0.142 -0.080 0.547 0.080 ;
      RECT 0.049 -0.080 0.142 0.260 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.316 1.120 0.900 1.280 ;
      RECT 0.224 0.909 0.316 1.280 ;
      RECT 0.000 1.120 0.224 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.049 0.742 0.491 0.796 ;
  END
END AOI211X1

MACRO AND3X1
  CLASS CORE ;
  FOREIGN AND3X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.796 0.274 0.859 0.989 ;
      RECT 0.734 0.274 0.796 0.355 ;
      RECT 0.758 0.829 0.796 0.989 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.397 0.408 0.539 0.511 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.184 0.677 0.322 0.786 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.426 0.158 0.548 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.638 -0.080 0.900 0.080 ;
      RECT 0.545 -0.080 0.638 0.122 ;
      RECT 0.000 -0.080 0.545 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.694 1.120 0.900 1.280 ;
      RECT 0.694 0.671 0.734 0.722 ;
      RECT 0.631 0.671 0.694 1.280 ;
      RECT 0.360 1.120 0.631 1.280 ;
      RECT 0.359 1.078 0.360 1.280 ;
      RECT 0.270 1.065 0.359 1.280 ;
      RECT 0.267 1.078 0.270 1.280 ;
      RECT 0.000 1.120 0.267 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.664 0.417 0.734 0.504 ;
      RECT 0.601 0.283 0.664 0.504 ;
      RECT 0.288 0.283 0.601 0.338 ;
      RECT 0.462 0.567 0.477 0.744 ;
      RECT 0.400 0.567 0.462 0.995 ;
      RECT 0.288 0.567 0.400 0.621 ;
      RECT 0.142 0.940 0.400 0.995 ;
      RECT 0.225 0.283 0.288 0.621 ;
      RECT 0.142 0.283 0.225 0.338 ;
      RECT 0.049 0.257 0.142 0.338 ;
      RECT 0.049 0.940 0.142 1.038 ;
  END
END AND3X1

MACRO AND2XL
  CLASS CORE ;
  FOREIGN AND2XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.624 0.567 0.663 0.633 ;
      RECT 0.563 0.344 0.624 0.845 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.219 0.564 0.320 0.702 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.040 0.433 0.150 0.551 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.475 -0.080 0.700 0.080 ;
      RECT 0.384 -0.080 0.475 0.122 ;
      RECT 0.000 -0.080 0.384 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.371 1.120 0.700 1.280 ;
      RECT 0.122 1.078 0.371 1.280 ;
      RECT 0.000 1.120 0.122 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.440 0.195 0.501 0.827 ;
      RECT 0.138 0.195 0.440 0.250 ;
      RECT 0.212 0.773 0.440 0.827 ;
      RECT 0.122 0.760 0.212 0.840 ;
      RECT 0.048 0.182 0.138 0.263 ;
  END
END AND2XL

MACRO AND2X4
  CLASS CORE ;
  FOREIGN AND2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.860 0.433 0.862 0.767 ;
      RECT 0.784 0.331 0.860 0.798 ;
      RECT 0.758 0.326 0.784 0.798 ;
      RECT 0.592 0.326 0.758 0.433 ;
      RECT 0.580 0.717 0.758 0.798 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.322 0.471 0.375 0.562 ;
      RECT 0.312 0.471 0.322 0.786 ;
      RECT 0.259 0.507 0.312 0.786 ;
      RECT 0.218 0.627 0.259 0.786 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.142 0.482 0.145 0.574 ;
      RECT 0.038 0.482 0.142 0.660 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.848 -0.080 0.900 0.080 ;
      RECT 0.755 -0.080 0.848 0.243 ;
      RECT 0.480 -0.080 0.755 0.080 ;
      RECT 0.387 -0.080 0.480 0.122 ;
      RECT 0.000 -0.080 0.387 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.848 1.120 0.900 1.280 ;
      RECT 0.755 0.914 0.848 1.280 ;
      RECT 0.487 1.120 0.755 1.280 ;
      RECT 0.394 1.078 0.487 1.280 ;
      RECT 0.146 1.120 0.394 1.280 ;
      RECT 0.046 1.078 0.146 1.280 ;
      RECT 0.000 1.120 0.046 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.503 0.498 0.663 0.579 ;
      RECT 0.449 0.354 0.503 0.671 ;
      RECT 0.440 0.354 0.449 0.910 ;
      RECT 0.142 0.354 0.440 0.408 ;
      RECT 0.386 0.617 0.440 0.910 ;
      RECT 0.202 0.855 0.386 0.910 ;
      RECT 0.049 0.343 0.142 0.424 ;
  END
END AND2X4

MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.642 0.227 0.654 0.767 ;
      RECT 0.593 0.195 0.642 1.002 ;
      RECT 0.582 0.195 0.593 0.439 ;
      RECT 0.552 0.688 0.593 1.002 ;
      RECT 0.552 0.195 0.582 0.390 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.833 0.361 0.935 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.138 0.504 0.202 0.585 ;
      RECT 0.037 0.504 0.138 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.440 -0.080 0.700 0.080 ;
      RECT 0.350 -0.080 0.440 0.122 ;
      RECT 0.000 -0.080 0.350 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.151 1.120 0.700 1.280 ;
      RECT 0.048 1.078 0.151 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.325 0.512 0.521 0.594 ;
      RECT 0.264 0.348 0.325 0.737 ;
      RECT 0.138 0.348 0.264 0.402 ;
      RECT 0.216 0.654 0.264 0.737 ;
      RECT 0.048 0.321 0.138 0.402 ;
  END
END AND2X2

MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.624 0.567 0.663 0.633 ;
      RECT 0.624 0.320 0.639 0.439 ;
      RECT 0.624 0.732 0.639 0.927 ;
      RECT 0.563 0.320 0.624 0.927 ;
      RECT 0.562 0.320 0.563 0.439 ;
      RECT 0.549 0.732 0.563 0.927 ;
      RECT 0.549 0.320 0.562 0.401 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.551 0.322 0.689 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.040 0.433 0.150 0.551 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.475 -0.080 0.700 0.080 ;
      RECT 0.384 -0.080 0.475 0.122 ;
      RECT 0.000 -0.080 0.384 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.465 1.120 0.700 1.280 ;
      RECT 0.347 1.078 0.465 1.280 ;
      RECT 0.209 1.120 0.347 1.280 ;
      RECT 0.119 1.078 0.209 1.280 ;
      RECT 0.000 1.120 0.119 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.487 0.461 0.500 0.561 ;
      RECT 0.426 0.195 0.487 0.827 ;
      RECT 0.138 0.195 0.426 0.250 ;
      RECT 0.423 0.461 0.426 0.561 ;
      RECT 0.209 0.773 0.426 0.827 ;
      RECT 0.119 0.760 0.209 0.840 ;
      RECT 0.048 0.182 0.138 0.263 ;
  END
END AND2X1

MACRO ADDHXL
  CLASS CORE ;
  FOREIGN ADDHXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.200 0.706 1.213 0.763 ;
      RECT 1.136 0.387 1.200 0.763 ;
      RECT 0.961 0.387 1.136 0.442 ;
      RECT 0.939 0.708 1.136 0.763 ;
      RECT 0.898 0.261 0.961 0.442 ;
      RECT 0.876 0.708 0.939 0.877 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.935 0.439 1.941 0.494 ;
      RECT 1.872 0.150 1.935 0.915 ;
      RECT 1.791 0.861 1.872 0.915 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.813 0.936 1.583 0.990 ;
      RECT 0.993 0.508 1.056 0.652 ;
      RECT 0.813 0.598 0.993 0.652 ;
      RECT 0.749 0.598 0.813 0.990 ;
      RECT 0.584 0.682 0.749 0.767 ;
      RECT 0.489 0.682 0.584 0.737 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.427 0.550 1.598 0.650 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.752 -0.080 2.000 0.080 ;
      RECT 1.658 -0.080 1.752 0.216 ;
      RECT 1.395 -0.080 1.658 0.080 ;
      RECT 1.302 -0.080 1.395 0.122 ;
      RECT 0.353 -0.080 1.302 0.080 ;
      RECT 0.259 -0.080 0.353 0.122 ;
      RECT 0.000 -0.080 0.259 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.729 1.120 2.000 1.280 ;
      RECT 1.635 1.078 1.729 1.280 ;
      RECT 1.307 1.120 1.635 1.280 ;
      RECT 1.213 1.078 1.307 1.280 ;
      RECT 0.353 1.120 1.213 1.280 ;
      RECT 0.259 1.078 0.353 1.280 ;
      RECT 0.000 1.120 0.259 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.736 0.669 1.802 0.765 ;
      RECT 1.672 0.331 1.736 0.765 ;
      RECT 1.621 0.331 1.672 0.386 ;
      RECT 1.501 0.711 1.672 0.765 ;
      RECT 1.438 0.711 1.501 0.877 ;
      RECT 1.298 0.275 1.361 0.877 ;
      RECT 1.160 0.275 1.298 0.330 ;
      RECT 1.059 0.823 1.298 0.877 ;
      RECT 1.096 0.150 1.160 0.330 ;
      RECT 0.825 0.150 1.096 0.205 ;
      RECT 0.762 0.150 0.825 0.508 ;
      RECT 0.383 0.454 0.762 0.508 ;
      RECT 0.634 0.151 0.697 0.246 ;
      RECT 0.621 0.852 0.685 1.008 ;
      RECT 0.255 0.301 0.668 0.356 ;
      RECT 0.128 0.192 0.634 0.246 ;
      RECT 0.128 0.954 0.621 1.008 ;
      RECT 0.423 0.844 0.507 0.899 ;
      RECT 0.360 0.711 0.423 0.899 ;
      RECT 0.320 0.454 0.383 0.636 ;
      RECT 0.255 0.711 0.360 0.765 ;
      RECT 0.191 0.301 0.255 0.765 ;
      RECT 0.065 0.192 0.128 1.008 ;
  END
END ADDHXL

MACRO ADDHX4
  CLASS CORE ;
  FOREIGN ADDHX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.742 0.158 2.824 0.239 ;
      RECT 2.157 0.158 2.742 0.213 ;
      RECT 1.518 0.711 2.716 0.765 ;
      RECT 2.096 0.158 2.157 0.392 ;
      RECT 2.043 0.300 2.096 0.392 ;
      RECT 1.538 0.337 2.043 0.392 ;
      RECT 1.518 0.300 1.538 0.633 ;
      RECT 1.457 0.300 1.518 0.765 ;
      RECT 1.437 0.300 1.457 0.633 ;
      RECT 1.267 0.711 1.457 0.765 ;
      RECT 1.384 0.313 1.437 0.405 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.648 0.567 4.688 0.900 ;
      RECT 4.587 0.338 4.648 0.900 ;
      RECT 4.537 0.338 4.587 0.393 ;
      RECT 4.416 0.665 4.587 0.720 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.238 0.463 2.640 0.518 ;
      RECT 2.234 0.463 2.238 0.618 ;
      RECT 2.173 0.463 2.234 0.627 ;
      RECT 2.157 0.563 2.173 0.627 ;
      RECT 1.694 0.563 2.157 0.618 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.288 0.488 4.111 0.543 ;
      RECT 3.227 0.439 3.288 0.543 ;
      RECT 3.207 0.439 3.227 0.494 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.797 -0.080 4.900 0.080 ;
      RECT 4.706 -0.080 4.797 0.214 ;
      RECT 4.457 -0.080 4.706 0.080 ;
      RECT 4.367 -0.080 4.457 0.214 ;
      RECT 4.101 -0.080 4.367 0.080 ;
      RECT 4.010 -0.080 4.101 0.211 ;
      RECT 3.761 -0.080 4.010 0.080 ;
      RECT 3.671 -0.080 3.761 0.211 ;
      RECT 3.422 -0.080 3.671 0.080 ;
      RECT 3.332 -0.080 3.422 0.198 ;
      RECT 1.241 -0.080 3.332 0.080 ;
      RECT 1.151 -0.080 1.241 0.122 ;
      RECT 0.827 -0.080 1.151 0.080 ;
      RECT 0.737 -0.080 0.827 0.122 ;
      RECT 0.477 -0.080 0.737 0.080 ;
      RECT 0.387 -0.080 0.477 0.214 ;
      RECT 0.138 -0.080 0.387 0.080 ;
      RECT 0.048 -0.080 0.138 0.211 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.705 1.120 4.900 1.280 ;
      RECT 4.586 1.078 4.705 1.280 ;
      RECT 4.331 1.120 4.586 1.280 ;
      RECT 4.241 0.989 4.331 1.280 ;
      RECT 3.985 1.120 4.241 1.280 ;
      RECT 3.895 0.989 3.985 1.280 ;
      RECT 3.646 1.120 3.895 1.280 ;
      RECT 3.556 0.989 3.646 1.280 ;
      RECT 3.295 1.120 3.556 1.280 ;
      RECT 3.204 1.078 3.295 1.280 ;
      RECT 2.881 1.120 3.204 1.280 ;
      RECT 2.791 1.078 2.881 1.280 ;
      RECT 1.188 1.120 2.791 1.280 ;
      RECT 1.098 1.078 1.188 1.280 ;
      RECT 0.827 1.120 1.098 1.280 ;
      RECT 0.737 1.078 0.827 1.280 ;
      RECT 0.477 1.120 0.737 1.280 ;
      RECT 0.387 0.989 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.989 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.285 0.499 4.443 0.554 ;
      RECT 4.224 0.499 4.285 0.658 ;
      RECT 3.577 0.355 4.270 0.410 ;
      RECT 3.086 0.604 4.224 0.658 ;
      RECT 3.261 0.715 4.156 0.770 ;
      RECT 3.501 0.324 3.577 0.410 ;
      RECT 3.243 0.324 3.501 0.379 ;
      RECT 3.200 0.715 3.261 0.876 ;
      RECT 3.182 0.170 3.243 0.379 ;
      RECT 2.838 0.821 3.200 0.876 ;
      RECT 2.946 0.170 3.182 0.225 ;
      RECT 3.068 0.604 3.086 0.744 ;
      RECT 3.007 0.331 3.068 0.744 ;
      RECT 2.992 0.689 3.007 0.744 ;
      RECT 2.885 0.170 2.946 0.392 ;
      RECT 2.838 0.337 2.885 0.392 ;
      RECT 2.777 0.337 2.838 1.004 ;
      RECT 2.239 0.337 2.777 0.392 ;
      RECT 2.127 0.949 2.777 1.004 ;
      RECT 2.066 0.876 2.127 1.004 ;
      RECT 1.428 0.876 2.066 0.931 ;
      RECT 1.368 0.158 1.969 0.213 ;
      RECT 1.310 0.987 1.867 1.042 ;
      RECT 1.367 0.842 1.428 0.931 ;
      RECT 1.307 0.158 1.368 0.248 ;
      RECT 0.770 0.842 1.367 0.896 ;
      RECT 0.993 0.361 1.319 0.415 ;
      RECT 1.249 0.954 1.310 1.042 ;
      RECT 0.762 0.193 1.307 0.248 ;
      RECT 0.647 0.954 1.249 1.008 ;
      RECT 0.932 0.361 0.993 0.733 ;
      RECT 0.711 0.519 0.770 0.896 ;
      RECT 0.701 0.193 0.762 0.392 ;
      RECT 0.709 0.493 0.711 0.896 ;
      RECT 0.247 0.493 0.709 0.574 ;
      RECT 0.184 0.337 0.701 0.392 ;
      RECT 0.586 0.665 0.647 1.008 ;
      RECT 0.184 0.665 0.586 0.720 ;
      RECT 0.123 0.337 0.184 0.720 ;
  END
END ADDHX4

MACRO ADDHX2
  CLASS CORE ;
  FOREIGN ADDHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.539 0.306 1.601 0.392 ;
      RECT 1.142 0.674 1.578 0.755 ;
      RECT 0.947 0.319 1.539 0.374 ;
      RECT 1.009 0.687 1.142 0.755 ;
      RECT 0.879 0.687 1.009 0.761 ;
      RECT 0.894 0.306 0.947 0.374 ;
      RECT 0.879 0.306 0.894 0.387 ;
      RECT 0.818 0.306 0.879 0.761 ;
      RECT 0.803 0.306 0.818 0.387 ;
      RECT 0.812 0.669 0.818 0.761 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.985 0.324 3.099 0.405 ;
      RECT 2.964 0.324 2.985 0.439 ;
      RECT 2.967 0.626 2.982 0.733 ;
      RECT 2.964 0.626 2.967 0.761 ;
      RECT 2.902 0.350 2.964 0.761 ;
      RECT 2.890 0.626 2.902 0.733 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.386 0.438 1.477 0.519 ;
      RECT 1.364 0.438 1.386 0.506 ;
      RECT 1.302 0.439 1.364 0.506 ;
      RECT 1.104 0.451 1.302 0.506 ;
      RECT 1.042 0.451 1.104 0.619 ;
      RECT 1.013 0.538 1.042 0.619 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.253 0.454 2.525 0.535 ;
      RECT 2.191 0.439 2.253 0.535 ;
      RECT 2.054 0.454 2.191 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.905 -0.080 3.200 0.080 ;
      RECT 2.813 -0.080 2.905 0.211 ;
      RECT 2.566 -0.080 2.813 0.080 ;
      RECT 2.474 -0.080 2.566 0.220 ;
      RECT 2.221 -0.080 2.474 0.080 ;
      RECT 2.129 -0.080 2.221 0.220 ;
      RECT 0.496 -0.080 2.129 0.080 ;
      RECT 0.404 -0.080 0.496 0.122 ;
      RECT 0.140 -0.080 0.404 0.080 ;
      RECT 0.048 -0.080 0.140 0.215 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.809 1.120 3.200 1.280 ;
      RECT 2.718 0.989 2.809 1.280 ;
      RECT 2.448 1.120 2.718 1.280 ;
      RECT 2.357 0.989 2.448 1.280 ;
      RECT 2.104 1.120 2.357 1.280 ;
      RECT 2.012 1.002 2.104 1.280 ;
      RECT 1.767 1.120 2.012 1.280 ;
      RECT 1.675 1.065 1.767 1.280 ;
      RECT 0.496 1.120 1.675 1.280 ;
      RECT 0.404 1.078 0.496 1.280 ;
      RECT 0.140 1.120 0.404 1.280 ;
      RECT 0.048 1.002 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.760 0.514 2.789 0.595 ;
      RECT 2.698 0.514 2.760 0.658 ;
      RECT 2.646 0.313 2.738 0.394 ;
      RECT 1.918 0.604 2.698 0.658 ;
      RECT 1.996 0.324 2.646 0.379 ;
      RECT 2.246 0.713 2.621 0.794 ;
      RECT 2.185 0.713 2.246 0.896 ;
      RECT 1.725 0.842 2.185 0.896 ;
      RECT 1.934 0.158 1.996 0.379 ;
      RECT 1.725 0.158 1.934 0.213 ;
      RECT 1.851 0.604 1.918 0.762 ;
      RECT 1.826 0.289 1.851 0.762 ;
      RECT 1.789 0.289 1.826 0.658 ;
      RECT 1.663 0.158 1.725 0.896 ;
      RECT 1.352 0.158 1.663 0.213 ;
      RECT 1.538 0.842 1.663 0.896 ;
      RECT 1.476 0.842 1.538 1.024 ;
      RECT 1.406 0.969 1.476 1.024 ;
      RECT 1.314 0.969 1.406 1.050 ;
      RECT 0.637 0.995 1.314 1.050 ;
      RECT 0.620 0.158 1.067 0.213 ;
      RECT 0.793 0.885 1.061 0.939 ;
      RECT 0.731 0.843 0.793 0.939 ;
      RECT 0.675 0.302 0.737 0.733 ;
      RECT 0.388 0.843 0.731 0.898 ;
      RECT 0.609 0.302 0.675 0.357 ;
      RECT 0.609 0.652 0.675 0.733 ;
      RECT 0.575 0.952 0.637 1.050 ;
      RECT 0.558 0.158 0.620 0.248 ;
      RECT 0.264 0.952 0.575 1.007 ;
      RECT 0.388 0.193 0.558 0.248 ;
      RECT 0.326 0.193 0.388 0.898 ;
      RECT 0.221 0.325 0.326 0.406 ;
      RECT 0.221 0.652 0.326 0.733 ;
      RECT 0.202 0.850 0.264 1.007 ;
      RECT 0.156 0.505 0.248 0.586 ;
      RECT 0.133 0.850 0.202 0.905 ;
      RECT 0.133 0.531 0.156 0.586 ;
      RECT 0.071 0.531 0.133 0.905 ;
  END
END ADDHX2

MACRO ADDHX1
  CLASS CORE ;
  FOREIGN ADDHX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.062 0.317 1.123 0.767 ;
      RECT 0.952 0.317 1.062 0.371 ;
      RECT 0.860 0.676 1.062 0.767 ;
      RECT 0.891 0.288 0.952 0.371 ;
      RECT 0.799 0.676 0.860 0.888 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.018 0.439 2.043 0.494 ;
      RECT 1.962 0.329 2.018 0.494 ;
      RECT 1.957 0.329 1.962 0.742 ;
      RECT 1.901 0.439 1.957 0.742 ;
      RECT 1.863 0.687 1.901 0.742 ;
      RECT 1.802 0.687 1.863 0.945 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.547 0.600 1.608 0.820 ;
      RECT 1.368 0.765 1.547 0.820 ;
      RECT 1.307 0.765 1.368 1.008 ;
      RECT 0.738 0.954 1.307 1.008 ;
      RECT 0.940 0.429 1.001 0.600 ;
      RECT 0.738 0.545 0.940 0.600 ;
      RECT 0.677 0.545 0.738 1.008 ;
      RECT 0.582 0.545 0.677 0.633 ;
      RECT 0.561 0.545 0.582 0.613 ;
      RECT 0.471 0.532 0.561 0.613 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.184 0.433 1.346 0.533 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.896 -0.080 2.100 0.080 ;
      RECT 1.835 -0.080 1.896 0.333 ;
      RECT 1.359 -0.080 1.835 0.080 ;
      RECT 1.807 0.283 1.835 0.333 ;
      RECT 1.746 0.283 1.807 0.395 ;
      RECT 1.269 -0.080 1.359 0.122 ;
      RECT 0.361 -0.080 1.269 0.080 ;
      RECT 0.270 -0.080 0.361 0.122 ;
      RECT 0.000 -0.080 0.270 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.718 1.120 2.100 1.280 ;
      RECT 1.628 1.078 1.718 1.280 ;
      RECT 1.267 1.120 1.628 1.280 ;
      RECT 1.177 1.078 1.267 1.280 ;
      RECT 0.339 1.120 1.177 1.280 ;
      RECT 0.249 1.078 0.339 1.280 ;
      RECT 0.000 1.120 0.249 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.730 0.471 1.814 0.552 ;
      RECT 1.684 0.158 1.774 0.213 ;
      RECT 1.684 0.471 1.730 0.930 ;
      RECT 1.669 0.158 1.684 0.930 ;
      RECT 1.623 0.158 1.669 0.526 ;
      RECT 1.491 0.875 1.669 0.930 ;
      RECT 1.485 0.288 1.560 0.369 ;
      RECT 1.430 0.875 1.491 0.962 ;
      RECT 1.470 0.288 1.485 0.711 ;
      RECT 1.424 0.301 1.470 0.711 ;
      RECT 1.246 0.301 1.424 0.356 ;
      RECT 1.246 0.656 1.424 0.711 ;
      RECT 1.185 0.192 1.246 0.356 ;
      RECT 1.185 0.656 1.246 0.899 ;
      RECT 1.157 0.192 1.185 0.246 ;
      RECT 0.976 0.844 1.185 0.899 ;
      RECT 1.067 0.161 1.157 0.246 ;
      RECT 0.830 0.161 1.067 0.215 ;
      RECT 0.769 0.161 0.830 0.465 ;
      RECT 0.367 0.411 0.769 0.465 ;
      RECT 0.647 0.150 0.708 0.246 ;
      RECT 0.245 0.301 0.676 0.356 ;
      RECT 0.123 0.192 0.647 0.246 ;
      RECT 0.555 0.954 0.616 1.049 ;
      RECT 0.123 0.954 0.555 1.008 ;
      RECT 0.398 0.757 0.488 0.838 ;
      RECT 0.245 0.757 0.398 0.812 ;
      RECT 0.306 0.411 0.367 0.610 ;
      RECT 0.184 0.301 0.245 0.812 ;
      RECT 0.062 0.181 0.123 1.008 ;
  END
END ADDHX1

MACRO ADDFX2
  CLASS CORE ;
  FOREIGN ADDFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.557 0.306 3.569 0.424 ;
      RECT 3.557 0.665 3.565 0.746 ;
      RECT 3.496 0.306 3.557 0.746 ;
      RECT 3.478 0.306 3.496 0.424 ;
      RECT 3.474 0.665 3.496 0.746 ;
      RECT 3.405 0.306 3.478 0.361 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.139 0.340 3.205 0.421 ;
      RECT 3.139 0.665 3.199 0.746 ;
      RECT 3.078 0.340 3.139 0.746 ;
      RECT 3.053 0.573 3.078 0.627 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.461 0.433 2.532 0.488 ;
      RECT 2.400 0.433 2.461 0.767 ;
      RECT 2.296 0.682 2.400 0.767 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.119 0.486 0.203 0.567 ;
      RECT 0.112 0.486 0.119 0.627 ;
      RECT 0.057 0.512 0.112 0.627 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.040 0.560 1.291 0.640 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.388 -0.080 3.700 0.080 ;
      RECT 3.297 -0.080 3.388 0.122 ;
      RECT 2.691 -0.080 3.297 0.080 ;
      RECT 2.600 -0.080 2.691 0.122 ;
      RECT 1.261 -0.080 2.600 0.080 ;
      RECT 1.171 -0.080 1.261 0.199 ;
      RECT 0.343 -0.080 1.171 0.080 ;
      RECT 0.252 -0.080 0.343 0.122 ;
      RECT 0.000 -0.080 0.252 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.384 1.120 3.700 1.280 ;
      RECT 3.293 1.078 3.384 1.280 ;
      RECT 2.385 1.120 3.293 1.280 ;
      RECT 2.294 1.078 2.385 1.280 ;
      RECT 0.320 1.120 2.294 1.280 ;
      RECT 0.230 1.078 0.320 1.280 ;
      RECT 0.000 1.120 0.230 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.373 0.480 3.434 0.569 ;
      RECT 3.341 0.514 3.373 0.569 ;
      RECT 3.280 0.514 3.341 0.939 ;
      RECT 2.791 0.885 3.280 0.939 ;
      RECT 2.508 0.995 3.034 1.050 ;
      RECT 2.971 0.150 3.013 0.205 ;
      RECT 2.971 0.743 2.983 0.824 ;
      RECT 2.910 0.150 2.971 0.824 ;
      RECT 2.535 0.193 2.910 0.248 ;
      RECT 2.892 0.743 2.910 0.824 ;
      RECT 2.790 0.320 2.848 0.562 ;
      RECT 2.790 0.765 2.791 0.939 ;
      RECT 2.787 0.320 2.790 0.939 ;
      RECT 2.730 0.507 2.787 0.939 ;
      RECT 2.728 0.507 2.730 0.846 ;
      RECT 2.700 0.765 2.728 0.846 ;
      RECT 2.595 0.302 2.656 0.685 ;
      RECT 2.412 0.302 2.595 0.357 ;
      RECT 2.584 0.630 2.595 0.685 ;
      RECT 2.523 0.630 2.584 0.846 ;
      RECT 2.473 0.150 2.535 0.248 ;
      RECT 2.447 0.954 2.508 1.050 ;
      RECT 1.570 0.150 2.473 0.205 ;
      RECT 2.097 0.954 2.447 1.008 ;
      RECT 2.351 0.260 2.412 0.357 ;
      RECT 1.781 0.260 2.351 0.314 ;
      RECT 2.288 0.523 2.339 0.604 ;
      RECT 2.226 0.377 2.288 0.604 ;
      RECT 2.220 0.549 2.226 0.604 ;
      RECT 2.158 0.549 2.220 0.898 ;
      RECT 2.096 0.852 2.097 1.008 ;
      RECT 2.036 0.377 2.096 1.008 ;
      RECT 2.034 0.377 2.036 0.907 ;
      RECT 1.915 0.852 2.034 0.907 ;
      RECT 1.911 0.426 1.973 0.798 ;
      RECT 1.903 0.426 1.911 0.481 ;
      RECT 1.814 0.743 1.911 0.798 ;
      RECT 1.842 0.377 1.903 0.481 ;
      RECT 1.781 0.562 1.850 0.643 ;
      RECT 1.785 0.743 1.814 0.915 ;
      RECT 1.753 0.743 1.785 1.050 ;
      RECT 1.719 0.260 1.781 0.688 ;
      RECT 1.723 0.835 1.753 1.050 ;
      RECT 1.403 0.965 1.723 1.050 ;
      RECT 1.648 0.632 1.719 0.688 ;
      RECT 1.415 0.493 1.658 0.576 ;
      RECT 1.622 0.632 1.648 0.815 ;
      RECT 1.587 0.632 1.622 0.829 ;
      RECT 1.539 0.748 1.587 0.829 ;
      RECT 1.508 0.150 1.570 0.417 ;
      RECT 1.531 0.748 1.539 0.911 ;
      RECT 1.478 0.761 1.531 0.911 ;
      RECT 1.479 0.270 1.508 0.417 ;
      RECT 1.109 0.270 1.479 0.325 ;
      RECT 0.918 0.856 1.478 0.911 ;
      RECT 1.353 0.389 1.415 0.801 ;
      RECT 0.443 0.995 1.403 1.050 ;
      RECT 0.986 0.389 1.353 0.444 ;
      RECT 1.041 0.746 1.353 0.801 ;
      RECT 1.048 0.208 1.109 0.325 ;
      RECT 0.654 0.208 1.048 0.263 ;
      RECT 0.980 0.710 1.041 0.801 ;
      RECT 0.925 0.343 0.986 0.444 ;
      RECT 0.857 0.721 0.918 0.911 ;
      RECT 0.849 0.721 0.857 0.776 ;
      RECT 0.788 0.494 0.849 0.776 ;
      RECT 0.734 0.832 0.796 0.940 ;
      RECT 0.777 0.494 0.788 0.549 ;
      RECT 0.715 0.338 0.777 0.549 ;
      RECT 0.567 0.832 0.734 0.887 ;
      RECT 0.654 0.604 0.699 0.752 ;
      RECT 0.638 0.208 0.654 0.752 ;
      RECT 0.593 0.208 0.638 0.658 ;
      RECT 0.531 0.726 0.567 0.887 ;
      RECT 0.506 0.332 0.531 0.887 ;
      RECT 0.470 0.332 0.506 0.781 ;
      RECT 0.402 0.700 0.470 0.781 ;
      RECT 0.382 0.870 0.443 1.050 ;
      RECT 0.368 0.486 0.398 0.567 ;
      RECT 0.330 0.870 0.382 0.925 ;
      RECT 0.330 0.332 0.368 0.567 ;
      RECT 0.307 0.332 0.330 0.925 ;
      RECT 0.139 0.332 0.307 0.387 ;
      RECT 0.268 0.499 0.307 0.925 ;
      RECT 0.048 0.688 0.268 0.769 ;
      RECT 0.048 0.194 0.139 0.387 ;
  END
END ADDFX2

MACRO ADDFX1
  CLASS CORE ;
  FOREIGN ADDFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.623 0.306 3.643 0.361 ;
      RECT 3.593 0.306 3.623 0.439 ;
      RECT 3.593 0.627 3.623 0.858 ;
      RECT 3.532 0.306 3.593 0.858 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.205 0.567 3.290 0.633 ;
      RECT 3.199 0.340 3.205 0.633 ;
      RECT 3.138 0.340 3.199 0.746 ;
      RECT 3.114 0.340 3.138 0.421 ;
      RECT 3.109 0.665 3.138 0.746 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.461 0.433 2.532 0.488 ;
      RECT 2.400 0.433 2.461 0.767 ;
      RECT 2.296 0.682 2.400 0.767 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.119 0.486 0.203 0.567 ;
      RECT 0.112 0.486 0.119 0.627 ;
      RECT 0.057 0.512 0.112 0.627 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.040 0.560 1.291 0.640 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.409 -0.080 3.700 0.080 ;
      RECT 3.318 -0.080 3.409 0.370 ;
      RECT 2.691 -0.080 3.318 0.080 ;
      RECT 2.600 -0.080 2.691 0.122 ;
      RECT 1.261 -0.080 2.600 0.080 ;
      RECT 1.171 -0.080 1.261 0.199 ;
      RECT 0.343 -0.080 1.171 0.080 ;
      RECT 0.252 -0.080 0.343 0.122 ;
      RECT 0.000 -0.080 0.252 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.410 1.120 3.700 1.280 ;
      RECT 3.320 0.951 3.410 1.280 ;
      RECT 2.385 1.120 3.320 1.280 ;
      RECT 2.294 1.078 2.385 1.280 ;
      RECT 0.320 1.120 2.294 1.280 ;
      RECT 0.230 1.078 0.320 1.280 ;
      RECT 0.000 1.120 0.230 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.373 0.480 3.434 0.856 ;
      RECT 3.109 0.801 3.373 0.856 ;
      RECT 3.047 0.801 3.109 0.939 ;
      RECT 2.508 0.995 3.058 1.050 ;
      RECT 2.791 0.885 3.047 0.939 ;
      RECT 2.974 0.150 3.015 0.205 ;
      RECT 2.974 0.743 2.983 0.824 ;
      RECT 2.912 0.150 2.974 0.824 ;
      RECT 2.910 0.150 2.912 0.248 ;
      RECT 2.892 0.743 2.912 0.824 ;
      RECT 2.535 0.193 2.910 0.248 ;
      RECT 2.791 0.320 2.851 0.421 ;
      RECT 2.790 0.320 2.791 0.939 ;
      RECT 2.730 0.367 2.790 0.939 ;
      RECT 2.700 0.765 2.730 0.846 ;
      RECT 2.597 0.302 2.659 0.685 ;
      RECT 2.412 0.302 2.597 0.357 ;
      RECT 2.584 0.630 2.597 0.685 ;
      RECT 2.523 0.630 2.584 0.846 ;
      RECT 2.473 0.150 2.535 0.248 ;
      RECT 2.447 0.954 2.508 1.050 ;
      RECT 1.570 0.150 2.473 0.205 ;
      RECT 2.097 0.954 2.447 1.008 ;
      RECT 2.351 0.260 2.412 0.357 ;
      RECT 1.781 0.260 2.351 0.314 ;
      RECT 2.288 0.523 2.339 0.604 ;
      RECT 2.226 0.377 2.288 0.604 ;
      RECT 2.220 0.549 2.226 0.604 ;
      RECT 2.158 0.549 2.220 0.898 ;
      RECT 2.096 0.852 2.097 1.008 ;
      RECT 2.036 0.377 2.096 1.008 ;
      RECT 2.034 0.377 2.036 0.907 ;
      RECT 1.915 0.852 2.034 0.907 ;
      RECT 1.911 0.426 1.973 0.798 ;
      RECT 1.903 0.426 1.911 0.481 ;
      RECT 1.814 0.743 1.911 0.798 ;
      RECT 1.842 0.377 1.903 0.481 ;
      RECT 1.781 0.562 1.850 0.643 ;
      RECT 1.785 0.743 1.814 0.900 ;
      RECT 1.753 0.743 1.785 1.050 ;
      RECT 1.719 0.260 1.781 0.688 ;
      RECT 1.723 0.819 1.753 1.050 ;
      RECT 1.403 0.965 1.723 1.050 ;
      RECT 1.648 0.632 1.719 0.688 ;
      RECT 1.415 0.493 1.658 0.576 ;
      RECT 1.622 0.632 1.648 0.815 ;
      RECT 1.587 0.632 1.622 0.829 ;
      RECT 1.539 0.748 1.587 0.829 ;
      RECT 1.508 0.150 1.570 0.417 ;
      RECT 1.531 0.748 1.539 0.911 ;
      RECT 1.478 0.761 1.531 0.911 ;
      RECT 1.479 0.270 1.508 0.417 ;
      RECT 1.109 0.270 1.479 0.325 ;
      RECT 0.918 0.856 1.478 0.911 ;
      RECT 1.353 0.389 1.415 0.801 ;
      RECT 0.443 0.995 1.403 1.050 ;
      RECT 0.986 0.389 1.353 0.444 ;
      RECT 1.041 0.746 1.353 0.801 ;
      RECT 1.048 0.208 1.109 0.325 ;
      RECT 0.654 0.208 1.048 0.263 ;
      RECT 0.980 0.710 1.041 0.801 ;
      RECT 0.925 0.343 0.986 0.444 ;
      RECT 0.857 0.721 0.918 0.911 ;
      RECT 0.849 0.721 0.857 0.776 ;
      RECT 0.788 0.494 0.849 0.776 ;
      RECT 0.734 0.832 0.796 0.940 ;
      RECT 0.777 0.494 0.788 0.549 ;
      RECT 0.715 0.338 0.777 0.549 ;
      RECT 0.567 0.832 0.734 0.887 ;
      RECT 0.654 0.604 0.699 0.777 ;
      RECT 0.638 0.208 0.654 0.777 ;
      RECT 0.593 0.208 0.638 0.658 ;
      RECT 0.531 0.726 0.567 0.887 ;
      RECT 0.506 0.332 0.531 0.887 ;
      RECT 0.470 0.332 0.506 0.781 ;
      RECT 0.402 0.700 0.470 0.781 ;
      RECT 0.382 0.870 0.443 1.050 ;
      RECT 0.368 0.486 0.398 0.567 ;
      RECT 0.330 0.870 0.382 0.925 ;
      RECT 0.330 0.332 0.368 0.567 ;
      RECT 0.307 0.332 0.330 0.925 ;
      RECT 0.139 0.332 0.307 0.387 ;
      RECT 0.268 0.499 0.307 0.925 ;
      RECT 0.048 0.688 0.268 0.769 ;
      RECT 0.048 0.194 0.139 0.387 ;
  END
END ADDFX1

MACRO ADDFHX4
  CLASS CORE ;
  FOREIGN ADDFHX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.849 0.433 5.889 0.767 ;
      RECT 5.788 0.333 5.849 0.767 ;
      RECT 5.733 0.333 5.788 0.414 ;
      RECT 5.733 0.671 5.788 0.752 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.501 0.433 5.540 0.767 ;
      RECT 5.440 0.346 5.501 0.767 ;
      RECT 5.395 0.346 5.440 0.401 ;
      RECT 5.394 0.671 5.440 0.752 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.016 0.567 5.192 0.658 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.603 0.635 3.715 0.715 ;
      RECT 3.542 0.635 3.603 0.761 ;
      RECT 3.377 0.635 3.542 0.715 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.191 0.433 0.329 0.571 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.992 -0.080 6.100 0.080 ;
      RECT 5.902 -0.080 5.992 0.233 ;
      RECT 5.654 -0.080 5.902 0.080 ;
      RECT 5.564 -0.080 5.654 0.233 ;
      RECT 5.295 -0.080 5.564 0.080 ;
      RECT 5.205 -0.080 5.295 0.122 ;
      RECT 3.586 -0.080 5.205 0.080 ;
      RECT 3.496 -0.080 3.586 0.122 ;
      RECT 0.864 -0.080 3.496 0.080 ;
      RECT 0.774 -0.080 0.864 0.122 ;
      RECT 0.330 -0.080 0.774 0.080 ;
      RECT 0.240 -0.080 0.330 0.122 ;
      RECT 0.000 -0.080 0.240 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.993 1.120 6.100 1.280 ;
      RECT 5.903 0.988 5.993 1.280 ;
      RECT 5.654 1.120 5.903 1.280 ;
      RECT 5.564 0.988 5.654 1.280 ;
      RECT 5.314 1.120 5.564 1.280 ;
      RECT 5.225 0.989 5.314 1.280 ;
      RECT 4.968 1.120 5.225 1.280 ;
      RECT 4.850 1.078 4.968 1.280 ;
      RECT 3.721 1.120 4.850 1.280 ;
      RECT 3.631 0.970 3.721 1.280 ;
      RECT 3.340 1.120 3.631 1.280 ;
      RECT 3.251 0.970 3.340 1.280 ;
      RECT 0.966 1.120 3.251 1.280 ;
      RECT 0.877 0.911 0.966 1.280 ;
      RECT 0.382 1.120 0.877 1.280 ;
      RECT 0.292 0.967 0.382 1.280 ;
      RECT 0.000 1.120 0.292 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.662 0.526 5.710 0.614 ;
      RECT 5.601 0.526 5.662 0.913 ;
      RECT 4.559 0.858 5.601 0.913 ;
      RECT 5.362 0.482 5.376 0.563 ;
      RECT 5.287 0.456 5.362 0.563 ;
      RECT 5.258 0.456 5.287 0.511 ;
      RECT 5.197 0.239 5.258 0.511 ;
      RECT 5.032 0.239 5.197 0.294 ;
      RECT 4.909 0.356 5.136 0.411 ;
      RECT 4.909 0.725 5.114 0.780 ;
      RECT 4.971 0.150 5.032 0.294 ;
      RECT 4.216 0.150 4.971 0.205 ;
      RECT 4.848 0.260 4.909 0.780 ;
      RECT 4.355 0.260 4.848 0.314 ;
      RECT 4.797 0.549 4.848 0.636 ;
      RECT 4.735 0.369 4.788 0.424 ;
      RECT 4.735 0.712 4.749 0.793 ;
      RECT 4.674 0.369 4.735 0.793 ;
      RECT 4.660 0.712 4.674 0.793 ;
      RECT 4.545 0.369 4.596 0.424 ;
      RECT 4.545 0.785 4.559 0.977 ;
      RECT 4.484 0.369 4.545 0.977 ;
      RECT 4.469 0.785 4.484 0.977 ;
      RECT 4.355 0.751 4.369 0.944 ;
      RECT 4.294 0.260 4.355 0.944 ;
      RECT 4.279 0.751 4.294 0.944 ;
      RECT 4.201 0.150 4.216 0.362 ;
      RECT 4.141 0.150 4.201 0.817 ;
      RECT 4.126 0.167 4.141 0.362 ;
      RECT 4.135 0.762 4.141 0.817 ;
      RECT 4.046 0.762 4.135 0.957 ;
      RECT 4.005 0.151 4.065 0.686 ;
      RECT 4.001 0.151 4.005 0.246 ;
      RECT 3.366 0.192 4.001 0.246 ;
      RECT 3.911 0.348 3.944 0.876 ;
      RECT 3.883 0.348 3.911 1.026 ;
      RECT 3.787 0.348 3.883 0.402 ;
      RECT 3.821 0.821 3.883 1.026 ;
      RECT 3.762 0.457 3.822 0.545 ;
      RECT 3.531 0.821 3.821 0.876 ;
      RECT 3.697 0.321 3.787 0.402 ;
      RECT 3.502 0.457 3.762 0.512 ;
      RECT 3.441 0.821 3.531 1.026 ;
      RECT 3.441 0.301 3.502 0.512 ;
      RECT 3.220 0.301 3.441 0.356 ;
      RECT 3.220 0.821 3.441 0.876 ;
      RECT 3.220 0.411 3.375 0.465 ;
      RECT 3.305 0.157 3.366 0.246 ;
      RECT 2.563 0.157 3.305 0.212 ;
      RECT 3.160 0.269 3.220 0.356 ;
      RECT 3.160 0.411 3.220 0.900 ;
      RECT 2.684 0.269 3.160 0.324 ;
      RECT 3.038 0.380 3.099 1.023 ;
      RECT 2.745 0.380 3.038 0.435 ;
      RECT 2.633 0.968 3.038 1.023 ;
      RECT 2.914 0.490 2.975 0.908 ;
      RECT 2.684 0.490 2.914 0.545 ;
      RECT 1.912 0.854 2.914 0.908 ;
      RECT 2.794 0.738 2.848 0.793 ;
      RECT 2.733 0.601 2.794 0.793 ;
      RECT 2.563 0.601 2.733 0.656 ;
      RECT 2.624 0.269 2.684 0.545 ;
      RECT 2.558 0.968 2.633 1.033 ;
      RECT 2.502 0.150 2.563 0.656 ;
      RECT 1.157 0.979 2.558 1.033 ;
      RECT 2.427 0.737 2.503 0.792 ;
      RECT 2.202 0.150 2.502 0.205 ;
      RECT 2.366 0.300 2.427 0.792 ;
      RECT 2.303 0.300 2.366 0.355 ;
      RECT 2.064 0.737 2.366 0.792 ;
      RECT 2.188 0.627 2.303 0.682 ;
      RECT 2.188 0.150 2.202 0.317 ;
      RECT 2.142 0.150 2.188 0.682 ;
      RECT 2.127 0.236 2.142 0.682 ;
      RECT 2.113 0.236 2.127 0.317 ;
      RECT 2.003 0.464 2.064 0.792 ;
      RECT 1.998 0.236 2.012 0.317 ;
      RECT 1.998 0.464 2.003 0.519 ;
      RECT 1.983 0.236 1.998 0.519 ;
      RECT 1.937 0.150 1.983 0.519 ;
      RECT 1.922 0.150 1.937 0.317 ;
      RECT 1.631 0.150 1.922 0.205 ;
      RECT 1.897 0.725 1.912 0.920 ;
      RECT 1.843 0.586 1.897 0.920 ;
      RECT 1.837 0.282 1.843 0.920 ;
      RECT 1.782 0.282 1.837 0.640 ;
      RECT 1.822 0.725 1.837 0.920 ;
      RECT 1.332 0.865 1.822 0.920 ;
      RECT 1.732 0.282 1.782 0.337 ;
      RECT 1.687 0.737 1.722 0.792 ;
      RECT 1.627 0.571 1.687 0.792 ;
      RECT 1.616 0.150 1.631 0.269 ;
      RECT 1.616 0.571 1.627 0.626 ;
      RECT 1.555 0.150 1.616 0.626 ;
      RECT 1.541 0.150 1.555 0.269 ;
      RECT 0.986 0.150 1.541 0.205 ;
      RECT 1.455 0.738 1.537 0.793 ;
      RECT 1.447 0.382 1.455 0.793 ;
      RECT 1.433 0.369 1.447 0.793 ;
      RECT 1.394 0.260 1.433 0.793 ;
      RECT 1.372 0.260 1.394 0.457 ;
      RECT 1.109 0.260 1.372 0.314 ;
      RECT 1.357 0.369 1.372 0.450 ;
      RECT 1.271 0.596 1.332 0.920 ;
      RECT 1.240 0.596 1.271 0.651 ;
      RECT 1.179 0.369 1.240 0.651 ;
      RECT 1.096 0.738 1.157 1.033 ;
      RECT 1.064 0.260 1.109 0.401 ;
      RECT 1.067 0.738 1.096 0.949 ;
      RECT 0.998 0.738 1.067 0.840 ;
      RECT 1.048 0.260 1.064 0.414 ;
      RECT 0.998 0.333 1.048 0.414 ;
      RECT 0.974 0.333 0.998 0.840 ;
      RECT 0.926 0.150 0.986 0.248 ;
      RECT 0.937 0.346 0.974 0.840 ;
      RECT 0.716 0.346 0.937 0.401 ;
      RECT 0.776 0.786 0.937 0.840 ;
      RECT 0.137 0.193 0.926 0.248 ;
      RECT 0.753 0.498 0.842 0.579 ;
      RECT 0.687 0.786 0.776 0.867 ;
      RECT 0.516 0.511 0.753 0.565 ;
      RECT 0.626 0.333 0.716 0.414 ;
      RECT 0.519 0.965 0.634 1.020 ;
      RECT 0.516 0.348 0.531 0.429 ;
      RECT 0.458 0.821 0.519 1.020 ;
      RECT 0.471 0.348 0.516 0.565 ;
      RECT 0.471 0.652 0.486 0.733 ;
      RECT 0.456 0.348 0.471 0.733 ;
      RECT 0.137 0.821 0.458 0.876 ;
      RECT 0.441 0.348 0.456 0.429 ;
      RECT 0.411 0.511 0.456 0.733 ;
      RECT 0.396 0.652 0.411 0.733 ;
      RECT 0.123 0.193 0.137 0.388 ;
      RECT 0.123 0.674 0.137 1.012 ;
      RECT 0.077 0.193 0.123 1.012 ;
      RECT 0.062 0.307 0.077 1.012 ;
      RECT 0.048 0.307 0.062 0.388 ;
      RECT 0.048 0.674 0.062 1.012 ;
  END
END ADDFHX4

MACRO ADDFHX2
  CLASS CORE ;
  FOREIGN ADDFHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.797 0.219 5.845 0.494 ;
      RECT 5.797 0.627 5.812 0.958 ;
      RECT 5.755 0.219 5.797 0.958 ;
      RECT 5.737 0.357 5.755 0.958 ;
      RECT 5.723 0.654 5.737 0.958 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.466 0.331 5.514 0.412 ;
      RECT 5.424 0.331 5.466 0.761 ;
      RECT 5.406 0.344 5.424 0.761 ;
      RECT 5.262 0.706 5.406 0.761 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.994 0.546 5.169 0.649 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.588 0.635 3.699 0.715 ;
      RECT 3.527 0.635 3.588 0.761 ;
      RECT 3.363 0.635 3.527 0.715 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.191 0.433 0.327 0.571 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.655 -0.080 5.900 0.080 ;
      RECT 5.566 -0.080 5.655 0.211 ;
      RECT 5.314 -0.080 5.566 0.080 ;
      RECT 5.224 -0.080 5.314 0.122 ;
      RECT 3.570 -0.080 5.224 0.080 ;
      RECT 3.481 -0.080 3.570 0.122 ;
      RECT 0.881 -0.080 3.481 0.080 ;
      RECT 0.791 -0.080 0.881 0.122 ;
      RECT 0.350 -0.080 0.791 0.080 ;
      RECT 0.260 -0.080 0.350 0.122 ;
      RECT 0.000 -0.080 0.260 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.623 1.120 5.900 1.280 ;
      RECT 5.533 0.988 5.623 1.280 ;
      RECT 5.291 1.120 5.533 1.280 ;
      RECT 5.202 0.988 5.291 1.280 ;
      RECT 4.940 1.120 5.202 1.280 ;
      RECT 4.834 1.078 4.940 1.280 ;
      RECT 3.705 1.120 4.834 1.280 ;
      RECT 3.615 0.970 3.705 1.280 ;
      RECT 3.326 1.120 3.615 1.280 ;
      RECT 3.237 0.970 3.326 1.280 ;
      RECT 0.962 1.120 3.237 1.280 ;
      RECT 0.873 0.911 0.962 1.280 ;
      RECT 0.380 1.120 0.873 1.280 ;
      RECT 0.291 0.967 0.380 1.280 ;
      RECT 0.000 1.120 0.291 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.527 0.526 5.587 0.913 ;
      RECT 4.539 0.858 5.527 0.913 ;
      RECT 5.278 0.239 5.339 0.579 ;
      RECT 5.010 0.239 5.278 0.294 ;
      RECT 4.888 0.356 5.114 0.411 ;
      RECT 4.888 0.744 5.092 0.799 ;
      RECT 4.950 0.150 5.010 0.294 ;
      RECT 4.183 0.150 4.950 0.205 ;
      RECT 4.827 0.260 4.888 0.799 ;
      RECT 4.336 0.260 4.827 0.314 ;
      RECT 4.776 0.549 4.827 0.636 ;
      RECT 4.714 0.369 4.767 0.424 ;
      RECT 4.714 0.721 4.729 0.802 ;
      RECT 4.654 0.369 4.714 0.802 ;
      RECT 4.639 0.721 4.654 0.802 ;
      RECT 4.525 0.369 4.576 0.424 ;
      RECT 4.525 0.785 4.539 0.977 ;
      RECT 4.464 0.369 4.525 0.977 ;
      RECT 4.450 0.785 4.464 0.977 ;
      RECT 4.336 0.751 4.350 0.944 ;
      RECT 4.275 0.260 4.336 0.944 ;
      RECT 4.261 0.751 4.275 0.944 ;
      RECT 4.123 0.150 4.183 0.798 ;
      RECT 4.117 0.743 4.123 0.798 ;
      RECT 4.042 0.743 4.117 0.975 ;
      RECT 3.987 0.151 4.048 0.686 ;
      RECT 4.028 0.780 4.042 0.975 ;
      RECT 3.983 0.151 3.987 0.246 ;
      RECT 3.351 0.192 3.983 0.246 ;
      RECT 3.879 0.335 3.927 0.726 ;
      RECT 3.879 0.819 3.894 1.014 ;
      RECT 3.866 0.335 3.879 1.014 ;
      RECT 3.770 0.335 3.866 0.389 ;
      RECT 3.819 0.671 3.866 1.014 ;
      RECT 3.805 0.819 3.819 1.014 ;
      RECT 3.745 0.457 3.806 0.545 ;
      RECT 3.515 0.824 3.805 0.879 ;
      RECT 3.681 0.321 3.770 0.402 ;
      RECT 3.486 0.457 3.745 0.512 ;
      RECT 3.426 0.824 3.515 1.025 ;
      RECT 3.426 0.301 3.486 0.512 ;
      RECT 3.206 0.301 3.426 0.356 ;
      RECT 3.206 0.824 3.426 0.879 ;
      RECT 3.206 0.411 3.360 0.465 ;
      RECT 3.290 0.157 3.351 0.246 ;
      RECT 2.552 0.157 3.290 0.212 ;
      RECT 3.146 0.269 3.206 0.356 ;
      RECT 3.146 0.411 3.206 0.900 ;
      RECT 2.673 0.269 3.146 0.324 ;
      RECT 3.025 0.380 3.085 1.023 ;
      RECT 2.733 0.380 3.025 0.435 ;
      RECT 2.621 0.968 3.025 1.023 ;
      RECT 2.901 0.490 2.962 0.910 ;
      RECT 2.673 0.490 2.901 0.545 ;
      RECT 1.889 0.855 2.901 0.910 ;
      RECT 2.782 0.738 2.836 0.793 ;
      RECT 2.721 0.601 2.782 0.793 ;
      RECT 2.552 0.601 2.721 0.656 ;
      RECT 2.612 0.269 2.673 0.545 ;
      RECT 2.546 0.968 2.621 1.050 ;
      RECT 2.491 0.150 2.552 0.656 ;
      RECT 1.156 0.995 2.546 1.050 ;
      RECT 2.416 0.737 2.493 0.792 ;
      RECT 2.178 0.150 2.491 0.205 ;
      RECT 2.356 0.300 2.416 0.792 ;
      RECT 2.293 0.300 2.356 0.355 ;
      RECT 2.011 0.737 2.356 0.792 ;
      RECT 2.178 0.627 2.293 0.682 ;
      RECT 2.118 0.150 2.178 0.682 ;
      RECT 1.989 0.293 2.011 0.792 ;
      RECT 1.951 0.150 1.989 0.792 ;
      RECT 1.929 0.150 1.951 0.348 ;
      RECT 1.609 0.150 1.929 0.205 ;
      RECT 1.829 0.446 1.889 0.919 ;
      RECT 1.800 0.446 1.829 0.501 ;
      RECT 1.326 0.864 1.829 0.919 ;
      RECT 1.739 0.269 1.800 0.501 ;
      RECT 1.685 0.724 1.714 0.805 ;
      RECT 1.625 0.571 1.685 0.805 ;
      RECT 1.609 0.571 1.625 0.626 ;
      RECT 1.549 0.150 1.609 0.626 ;
      RECT 1.003 0.150 1.549 0.205 ;
      RECT 1.470 0.725 1.530 0.806 ;
      RECT 1.441 0.260 1.470 0.806 ;
      RECT 1.409 0.260 1.441 0.793 ;
      RECT 1.125 0.260 1.409 0.314 ;
      RECT 1.387 0.369 1.409 0.457 ;
      RECT 1.266 0.596 1.326 0.919 ;
      RECT 1.255 0.596 1.266 0.651 ;
      RECT 1.195 0.369 1.255 0.651 ;
      RECT 1.095 0.785 1.156 1.050 ;
      RECT 1.065 0.260 1.125 0.370 ;
      RECT 1.058 0.785 1.095 0.852 ;
      RECT 0.994 0.315 1.065 0.370 ;
      RECT 0.994 0.785 1.058 0.839 ;
      RECT 0.943 0.150 1.003 0.248 ;
      RECT 0.933 0.315 0.994 0.839 ;
      RECT 0.137 0.193 0.943 0.248 ;
      RECT 0.734 0.315 0.933 0.370 ;
      RECT 0.776 0.785 0.933 0.839 ;
      RECT 0.770 0.498 0.860 0.579 ;
      RECT 0.678 0.785 0.776 0.852 ;
      RECT 0.535 0.511 0.770 0.565 ;
      RECT 0.644 0.302 0.734 0.383 ;
      RECT 0.517 0.965 0.631 1.020 ;
      RECT 0.535 0.348 0.550 0.429 ;
      RECT 0.484 0.348 0.535 0.565 ;
      RECT 0.456 0.821 0.517 1.020 ;
      RECT 0.475 0.348 0.484 0.733 ;
      RECT 0.460 0.348 0.475 0.429 ;
      RECT 0.423 0.511 0.475 0.733 ;
      RECT 0.137 0.821 0.456 0.876 ;
      RECT 0.394 0.652 0.423 0.733 ;
      RECT 0.122 0.193 0.137 0.369 ;
      RECT 0.122 0.674 0.137 1.012 ;
      RECT 0.076 0.193 0.122 1.012 ;
      RECT 0.062 0.288 0.076 1.012 ;
      RECT 0.047 0.288 0.062 0.369 ;
      RECT 0.047 0.674 0.062 1.012 ;
  END
END ADDFHX2

MACRO ADDFHX1
  CLASS CORE ;
  FOREIGN ADDFHX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.938 0.439 3.943 0.494 ;
      RECT 3.877 0.326 3.938 0.838 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.590 0.439 3.596 0.494 ;
      RECT 3.530 0.326 3.590 0.877 ;
      RECT 3.455 0.823 3.530 0.877 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.325 0.700 3.422 0.761 ;
      RECT 3.265 0.560 3.325 0.761 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.819 0.700 2.030 0.804 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.188 0.439 0.291 0.593 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.805 -0.080 4.000 0.080 ;
      RECT 3.715 -0.080 3.805 0.122 ;
      RECT 3.448 -0.080 3.715 0.080 ;
      RECT 3.358 -0.080 3.448 0.122 ;
      RECT 2.017 -0.080 3.358 0.080 ;
      RECT 1.928 -0.080 2.017 0.122 ;
      RECT 0.464 -0.080 1.928 0.080 ;
      RECT 0.374 -0.080 0.464 0.122 ;
      RECT 0.000 -0.080 0.374 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.744 1.120 4.000 1.280 ;
      RECT 3.655 1.078 3.744 1.280 ;
      RECT 3.157 1.120 3.655 1.280 ;
      RECT 3.067 1.078 3.157 1.280 ;
      RECT 1.972 1.120 3.067 1.280 ;
      RECT 1.883 0.983 1.972 1.280 ;
      RECT 0.628 1.120 1.883 1.280 ;
      RECT 0.539 0.894 0.628 1.280 ;
      RECT 0.327 1.120 0.539 1.280 ;
      RECT 0.237 0.909 0.327 1.280 ;
      RECT 0.000 1.120 0.237 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.746 0.585 3.769 0.670 ;
      RECT 3.685 0.585 3.746 1.008 ;
      RECT 2.752 0.954 3.685 1.008 ;
      RECT 3.298 0.192 3.634 0.246 ;
      RECT 3.177 0.357 3.403 0.412 ;
      RECT 3.177 0.824 3.358 0.879 ;
      RECT 3.237 0.150 3.298 0.246 ;
      RECT 2.486 0.150 3.237 0.205 ;
      RECT 3.116 0.260 3.177 0.879 ;
      RECT 2.661 0.260 3.116 0.314 ;
      RECT 3.028 0.610 3.116 0.664 ;
      RECT 3.024 0.386 3.055 0.440 ;
      RECT 2.967 0.386 3.024 0.551 ;
      RECT 2.963 0.386 2.967 0.879 ;
      RECT 2.906 0.496 2.963 0.879 ;
      RECT 2.867 0.824 2.906 0.879 ;
      RECT 2.833 0.386 2.866 0.440 ;
      RECT 2.772 0.386 2.833 0.765 ;
      RECT 2.752 0.711 2.772 0.765 ;
      RECT 2.692 0.711 2.752 1.008 ;
      RECT 2.601 0.260 2.661 0.655 ;
      RECT 2.563 0.600 2.601 0.655 ;
      RECT 2.502 0.600 2.563 0.893 ;
      RECT 2.441 0.150 2.486 0.440 ;
      RECT 2.426 0.150 2.441 1.023 ;
      RECT 2.381 0.386 2.426 1.023 ;
      RECT 2.262 0.968 2.381 1.023 ;
      RECT 2.161 0.152 2.347 0.207 ;
      RECT 2.260 0.373 2.320 0.913 ;
      RECT 2.221 0.373 2.260 0.454 ;
      RECT 2.177 0.858 2.260 0.913 ;
      RECT 2.161 0.586 2.199 0.780 ;
      RECT 2.063 0.858 2.177 0.951 ;
      RECT 2.138 0.152 2.161 0.780 ;
      RECT 2.100 0.152 2.138 0.640 ;
      RECT 1.867 0.206 2.100 0.261 ;
      RECT 1.768 0.858 2.063 0.913 ;
      RECT 1.979 0.324 2.040 0.620 ;
      RECT 1.746 0.324 1.979 0.379 ;
      RECT 1.806 0.150 1.867 0.261 ;
      RECT 1.382 0.150 1.806 0.205 ;
      RECT 1.747 0.858 1.768 0.982 ;
      RECT 1.686 0.496 1.747 0.982 ;
      RECT 1.685 0.260 1.746 0.379 ;
      RECT 1.503 0.260 1.685 0.314 ;
      RECT 1.564 0.369 1.625 1.049 ;
      RECT 0.813 0.994 1.564 1.049 ;
      RECT 1.443 0.260 1.503 0.939 ;
      RECT 1.003 0.885 1.443 0.939 ;
      RECT 1.321 0.150 1.382 0.805 ;
      RECT 1.132 0.179 1.192 0.805 ;
      RECT 0.586 0.179 1.132 0.233 ;
      RECT 1.003 0.290 1.017 0.371 ;
      RECT 0.942 0.290 1.003 0.939 ;
      RECT 0.928 0.290 0.942 0.371 ;
      RECT 0.813 0.290 0.827 0.371 ;
      RECT 0.752 0.290 0.813 1.049 ;
      RECT 0.738 0.290 0.752 0.371 ;
      RECT 0.560 0.480 0.686 0.573 ;
      RECT 0.526 0.179 0.586 0.261 ;
      RECT 0.499 0.361 0.560 0.769 ;
      RECT 0.123 0.206 0.526 0.261 ;
      RECT 0.406 0.361 0.499 0.415 ;
      RECT 0.395 0.714 0.499 0.769 ;
      RECT 0.123 0.723 0.137 0.946 ;
      RECT 0.062 0.206 0.123 0.946 ;
      RECT 0.047 0.723 0.062 0.946 ;
  END
END ADDFHX1

MACRO XOR3X4
  CLASS CORE ;
  FOREIGN XOR3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.977 0.700 4.990 1.033 ;
      RECT 4.964 0.227 4.977 1.033 ;
      RECT 4.916 0.199 4.964 1.033 ;
      RECT 4.874 0.199 4.916 0.392 ;
      RECT 4.890 0.652 4.916 1.033 ;
      RECT 4.885 0.652 4.890 0.733 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.557 0.936 4.646 1.017 ;
      RECT 4.450 0.962 4.557 1.017 ;
      RECT 4.390 0.962 4.450 1.027 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.152 0.637 3.180 0.718 ;
      RECT 3.091 0.375 3.152 0.718 ;
      RECT 3.025 0.375 3.091 0.500 ;
      RECT 3.003 0.439 3.025 0.500 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.290 0.526 0.386 0.607 ;
      RECT 0.230 0.526 0.290 0.627 ;
      RECT 0.173 0.526 0.230 0.607 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 -0.080 5.200 0.080 ;
      RECT 5.063 -0.080 5.153 0.377 ;
      RECT 4.764 -0.080 5.063 0.080 ;
      RECT 4.675 -0.080 4.764 0.135 ;
      RECT 2.462 -0.080 4.675 0.080 ;
      RECT 2.373 -0.080 2.462 0.122 ;
      RECT 2.010 -0.080 2.373 0.080 ;
      RECT 1.921 -0.080 2.010 0.122 ;
      RECT 1.601 -0.080 1.921 0.080 ;
      RECT 1.511 -0.080 1.601 0.122 ;
      RECT 0.336 -0.080 1.511 0.080 ;
      RECT 0.247 -0.080 0.336 0.359 ;
      RECT 0.000 -0.080 0.247 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 1.120 5.200 1.280 ;
      RECT 5.063 0.953 5.153 1.280 ;
      RECT 4.796 1.120 5.063 1.280 ;
      RECT 4.706 0.953 4.796 1.280 ;
      RECT 2.365 1.120 4.706 1.280 ;
      RECT 2.276 1.065 2.365 1.280 ;
      RECT 1.966 1.120 2.276 1.280 ;
      RECT 1.876 1.021 1.966 1.280 ;
      RECT 1.567 1.120 1.876 1.280 ;
      RECT 1.477 1.021 1.567 1.280 ;
      RECT 0.331 1.120 1.477 1.280 ;
      RECT 0.242 0.953 0.331 1.280 ;
      RECT 0.000 1.120 0.242 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.824 0.507 4.856 0.588 ;
      RECT 4.764 0.507 4.824 0.881 ;
      RECT 4.223 0.826 4.764 0.881 ;
      RECT 4.546 0.348 4.606 0.429 ;
      RECT 4.546 0.652 4.596 0.733 ;
      RECT 4.486 0.348 4.546 0.733 ;
      RECT 4.457 0.490 4.486 0.571 ;
      RECT 4.394 0.150 4.423 0.348 ;
      RECT 4.394 0.661 4.412 0.742 ;
      RECT 4.333 0.150 4.394 0.742 ;
      RECT 3.656 0.150 4.333 0.205 ;
      RECT 4.323 0.661 4.333 0.742 ;
      RECT 4.219 0.260 4.234 0.340 ;
      RECT 4.219 0.713 4.223 0.906 ;
      RECT 4.159 0.260 4.219 0.906 ;
      RECT 4.144 0.260 4.159 0.340 ;
      RECT 4.134 0.713 4.159 0.906 ;
      RECT 3.845 0.260 4.144 0.314 ;
      RECT 4.016 0.369 4.044 0.424 ;
      RECT 4.016 0.713 4.034 0.906 ;
      RECT 4.005 0.369 4.016 0.906 ;
      RECT 3.955 0.369 4.005 1.050 ;
      RECT 3.945 0.713 3.955 1.050 ;
      RECT 2.486 0.995 3.945 1.050 ;
      RECT 3.826 0.260 3.845 0.340 ;
      RECT 3.826 0.713 3.845 0.906 ;
      RECT 3.766 0.260 3.826 0.906 ;
      RECT 3.756 0.260 3.766 0.340 ;
      RECT 3.756 0.713 3.766 0.906 ;
      RECT 3.595 0.150 3.656 0.906 ;
      RECT 3.566 0.150 3.595 0.352 ;
      RECT 3.566 0.713 3.595 0.906 ;
      RECT 3.301 0.168 3.566 0.223 ;
      RECT 3.456 0.721 3.467 0.940 ;
      RECT 3.396 0.290 3.456 0.940 ;
      RECT 3.367 0.290 3.396 0.371 ;
      RECT 3.377 0.721 3.396 0.940 ;
      RECT 2.607 0.886 3.377 0.940 ;
      RECT 3.241 0.168 3.301 0.831 ;
      RECT 3.178 0.239 3.241 0.320 ;
      RECT 3.188 0.776 3.241 0.831 ;
      RECT 2.923 0.265 3.178 0.320 ;
      RECT 2.727 0.776 3.066 0.831 ;
      RECT 2.649 0.150 3.028 0.205 ;
      RECT 2.863 0.265 2.923 0.721 ;
      RECT 2.739 0.265 2.863 0.346 ;
      RECT 2.788 0.667 2.863 0.721 ;
      RECT 2.667 0.655 2.727 0.831 ;
      RECT 2.649 0.655 2.667 0.736 ;
      RECT 2.588 0.150 2.649 0.736 ;
      RECT 2.546 0.831 2.607 0.940 ;
      RECT 2.550 0.192 2.588 0.412 ;
      RECT 1.961 0.192 2.550 0.246 ;
      RECT 2.528 0.831 2.546 0.886 ;
      RECT 2.467 0.476 2.528 0.886 ;
      RECT 2.425 0.940 2.486 1.050 ;
      RECT 2.373 0.476 2.467 0.531 ;
      RECT 2.087 0.940 2.425 0.995 ;
      RECT 2.318 0.625 2.407 0.706 ;
      RECT 2.312 0.302 2.373 0.531 ;
      RECT 2.252 0.625 2.318 0.680 ;
      RECT 2.089 0.302 2.312 0.357 ;
      RECT 2.223 0.412 2.252 0.680 ;
      RECT 2.163 0.412 2.223 0.842 ;
      RECT 1.616 0.787 2.163 0.842 ;
      RECT 2.029 0.302 2.089 0.732 ;
      RECT 2.026 0.896 2.087 0.995 ;
      RECT 1.782 0.677 2.029 0.732 ;
      RECT 1.417 0.896 2.026 0.951 ;
      RECT 1.871 0.192 1.961 0.610 ;
      RECT 1.317 0.192 1.871 0.246 ;
      RECT 1.782 0.348 1.811 0.429 ;
      RECT 1.722 0.301 1.782 0.732 ;
      RECT 1.245 0.301 1.722 0.356 ;
      RECT 1.677 0.677 1.722 0.732 ;
      RECT 1.556 0.424 1.616 0.842 ;
      RECT 1.367 0.424 1.556 0.479 ;
      RECT 1.296 0.787 1.556 0.842 ;
      RECT 1.401 0.570 1.430 0.651 ;
      RECT 1.356 0.896 1.417 0.964 ;
      RECT 1.341 0.570 1.401 0.732 ;
      RECT 1.102 0.910 1.356 0.964 ;
      RECT 1.202 0.677 1.341 0.732 ;
      RECT 1.228 0.150 1.317 0.246 ;
      RECT 1.236 0.787 1.296 0.855 ;
      RECT 1.184 0.301 1.245 0.450 ;
      RECT 0.751 0.800 1.236 0.855 ;
      RECT 0.536 0.150 1.228 0.205 ;
      RECT 0.924 0.395 1.184 0.450 ;
      RECT 1.035 0.260 1.124 0.340 ;
      RECT 1.012 0.910 1.102 0.990 ;
      RECT 0.725 0.260 1.035 0.314 ;
      RECT 0.699 0.910 1.012 0.964 ;
      RECT 0.896 0.369 0.924 0.450 ;
      RECT 0.896 0.664 0.902 0.745 ;
      RECT 0.835 0.369 0.896 0.745 ;
      RECT 0.813 0.664 0.835 0.745 ;
      RECT 0.691 0.536 0.751 0.855 ;
      RECT 0.696 0.260 0.725 0.340 ;
      RECT 0.630 0.910 0.699 0.990 ;
      RECT 0.636 0.260 0.696 0.481 ;
      RECT 0.630 0.426 0.636 0.481 ;
      RECT 0.609 0.426 0.630 0.990 ;
      RECT 0.570 0.426 0.609 0.977 ;
      RECT 0.509 0.150 0.536 0.371 ;
      RECT 0.449 0.150 0.509 0.771 ;
      RECT 0.446 0.150 0.449 0.371 ;
      RECT 0.420 0.688 0.449 0.771 ;
      RECT 0.152 0.688 0.420 0.743 ;
      RECT 0.108 0.688 0.152 0.771 ;
      RECT 0.108 0.182 0.137 0.375 ;
      RECT 0.047 0.182 0.108 0.771 ;
  END
END XOR3X4

MACRO XOR3X2
  CLASS CORE ;
  FOREIGN XOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.152 0.227 3.165 0.720 ;
      RECT 3.142 0.199 3.152 0.733 ;
      RECT 3.103 0.199 3.142 0.761 ;
      RECT 3.060 0.199 3.103 0.392 ;
      RECT 3.080 0.652 3.103 0.761 ;
      RECT 3.060 0.652 3.080 0.733 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.672 0.788 2.815 0.900 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.892 0.573 1.898 0.627 ;
      RECT 1.863 0.573 1.892 0.769 ;
      RECT 1.801 0.426 1.863 0.769 ;
      RECT 1.714 0.426 1.801 0.507 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.120 0.526 0.221 0.607 ;
      RECT 0.058 0.526 0.120 0.627 ;
      RECT 0.038 0.526 0.058 0.607 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.947 -0.080 3.200 0.080 ;
      RECT 2.855 -0.080 2.947 0.135 ;
      RECT 0.995 -0.080 2.855 0.080 ;
      RECT 0.904 -0.080 0.995 0.179 ;
      RECT 0.140 -0.080 0.904 0.080 ;
      RECT 0.048 -0.080 0.140 0.359 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.968 1.120 3.200 1.280 ;
      RECT 2.877 0.953 2.968 1.280 ;
      RECT 0.952 1.120 2.877 1.280 ;
      RECT 0.861 1.011 0.952 1.280 ;
      RECT 0.162 1.120 0.861 1.280 ;
      RECT 0.070 0.953 0.162 1.280 ;
      RECT 0.000 1.120 0.070 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.998 0.507 3.041 0.588 ;
      RECT 2.936 0.238 2.998 0.588 ;
      RECT 2.742 0.238 2.936 0.293 ;
      RECT 2.723 0.348 2.785 0.429 ;
      RECT 2.723 0.652 2.774 0.733 ;
      RECT 2.680 0.182 2.742 0.293 ;
      RECT 2.661 0.348 2.723 0.733 ;
      RECT 2.392 0.182 2.680 0.237 ;
      RECT 2.632 0.490 2.661 0.571 ;
      RECT 2.567 0.292 2.597 0.373 ;
      RECT 2.567 0.713 2.586 0.906 ;
      RECT 2.556 0.292 2.567 0.906 ;
      RECT 2.505 0.292 2.556 1.050 ;
      RECT 2.494 0.713 2.505 1.050 ;
      RECT 1.243 0.995 2.494 1.050 ;
      RECT 2.373 0.150 2.392 0.343 ;
      RECT 2.373 0.713 2.392 0.906 ;
      RECT 2.311 0.150 2.373 0.906 ;
      RECT 2.300 0.150 2.311 0.343 ;
      RECT 2.300 0.713 2.311 0.906 ;
      RECT 2.136 0.150 2.198 0.906 ;
      RECT 2.106 0.150 2.136 0.352 ;
      RECT 2.106 0.713 2.136 0.906 ;
      RECT 1.653 0.150 2.106 0.205 ;
      RECT 1.982 0.290 2.044 0.940 ;
      RECT 1.902 0.290 1.982 0.371 ;
      RECT 1.912 0.860 1.982 0.940 ;
      RECT 1.367 0.886 1.912 0.940 ;
      RECT 1.647 0.655 1.739 0.736 ;
      RECT 1.623 0.150 1.653 0.412 ;
      RECT 1.623 0.655 1.647 0.710 ;
      RECT 1.591 0.150 1.623 0.710 ;
      RECT 1.561 0.219 1.591 0.710 ;
      RECT 1.491 0.776 1.545 0.831 ;
      RECT 1.459 0.249 1.491 0.831 ;
      RECT 1.429 0.200 1.459 0.831 ;
      RECT 1.367 0.200 1.429 0.304 ;
      RECT 0.871 0.249 1.367 0.304 ;
      RECT 1.305 0.358 1.367 0.940 ;
      RECT 0.995 0.358 1.305 0.413 ;
      RECT 1.230 0.468 1.243 0.523 ;
      RECT 1.181 0.887 1.243 1.050 ;
      RECT 1.200 0.468 1.230 0.667 ;
      RECT 1.138 0.468 1.200 0.832 ;
      RECT 0.539 0.887 1.181 0.942 ;
      RECT 0.593 0.777 1.138 0.832 ;
      RECT 0.933 0.358 0.995 0.723 ;
      RECT 0.718 0.668 0.933 0.723 ;
      RECT 0.842 0.249 0.871 0.610 ;
      RECT 0.780 0.150 0.842 0.610 ;
      RECT 0.345 0.150 0.780 0.205 ;
      RECT 0.656 0.267 0.718 0.723 ;
      RECT 0.531 0.493 0.593 0.832 ;
      RECT 0.469 0.260 0.539 0.340 ;
      RECT 0.469 0.887 0.539 0.968 ;
      RECT 0.447 0.260 0.469 0.968 ;
      RECT 0.407 0.273 0.447 0.955 ;
      RECT 0.283 0.150 0.345 0.745 ;
      RECT 0.253 0.150 0.283 0.350 ;
      RECT 0.253 0.664 0.283 0.745 ;
  END
END XOR3X2

MACRO XNOR3X4
  CLASS CORE ;
  FOREIGN XNOR3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.977 0.700 4.990 1.033 ;
      RECT 4.964 0.227 4.977 1.033 ;
      RECT 4.916 0.199 4.964 1.033 ;
      RECT 4.874 0.199 4.916 0.392 ;
      RECT 4.890 0.652 4.916 1.033 ;
      RECT 4.885 0.652 4.890 0.733 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.557 0.936 4.646 1.017 ;
      RECT 4.450 0.962 4.557 1.017 ;
      RECT 4.390 0.962 4.450 1.027 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.141 0.637 3.170 0.718 ;
      RECT 3.081 0.375 3.141 0.718 ;
      RECT 3.025 0.375 3.081 0.500 ;
      RECT 3.003 0.439 3.025 0.500 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.290 0.526 0.386 0.607 ;
      RECT 0.230 0.526 0.290 0.627 ;
      RECT 0.173 0.526 0.230 0.607 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 -0.080 5.200 0.080 ;
      RECT 5.063 -0.080 5.153 0.377 ;
      RECT 4.764 -0.080 5.063 0.080 ;
      RECT 4.675 -0.080 4.764 0.135 ;
      RECT 2.462 -0.080 4.675 0.080 ;
      RECT 2.373 -0.080 2.462 0.122 ;
      RECT 2.010 -0.080 2.373 0.080 ;
      RECT 1.921 -0.080 2.010 0.122 ;
      RECT 1.601 -0.080 1.921 0.080 ;
      RECT 1.511 -0.080 1.601 0.122 ;
      RECT 0.336 -0.080 1.511 0.080 ;
      RECT 0.247 -0.080 0.336 0.359 ;
      RECT 0.000 -0.080 0.247 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 1.120 5.200 1.280 ;
      RECT 5.063 0.953 5.153 1.280 ;
      RECT 4.796 1.120 5.063 1.280 ;
      RECT 4.706 0.953 4.796 1.280 ;
      RECT 2.365 1.120 4.706 1.280 ;
      RECT 2.276 1.065 2.365 1.280 ;
      RECT 1.966 1.120 2.276 1.280 ;
      RECT 1.876 1.021 1.966 1.280 ;
      RECT 1.567 1.120 1.876 1.280 ;
      RECT 1.477 1.021 1.567 1.280 ;
      RECT 0.331 1.120 1.477 1.280 ;
      RECT 0.242 0.953 0.331 1.280 ;
      RECT 0.000 1.120 0.242 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.824 0.507 4.856 0.588 ;
      RECT 4.764 0.507 4.824 0.881 ;
      RECT 4.230 0.826 4.764 0.881 ;
      RECT 4.554 0.348 4.617 0.429 ;
      RECT 4.554 0.652 4.596 0.733 ;
      RECT 4.494 0.348 4.554 0.733 ;
      RECT 4.457 0.499 4.494 0.580 ;
      RECT 4.394 0.348 4.433 0.429 ;
      RECT 4.394 0.661 4.412 0.742 ;
      RECT 4.333 0.150 4.394 0.742 ;
      RECT 3.645 0.150 4.333 0.205 ;
      RECT 4.323 0.661 4.333 0.742 ;
      RECT 4.230 0.260 4.244 0.352 ;
      RECT 4.223 0.260 4.230 0.881 ;
      RECT 4.169 0.260 4.223 0.906 ;
      RECT 4.155 0.260 4.169 0.352 ;
      RECT 4.134 0.713 4.169 0.906 ;
      RECT 3.834 0.260 4.155 0.314 ;
      RECT 4.016 0.369 4.044 0.424 ;
      RECT 4.016 0.713 4.034 0.906 ;
      RECT 4.005 0.369 4.016 0.906 ;
      RECT 3.955 0.369 4.005 1.050 ;
      RECT 3.945 0.713 3.955 1.050 ;
      RECT 2.486 0.995 3.945 1.050 ;
      RECT 3.826 0.713 3.845 0.906 ;
      RECT 3.826 0.260 3.834 0.352 ;
      RECT 3.766 0.260 3.826 0.906 ;
      RECT 3.745 0.260 3.766 0.352 ;
      RECT 3.756 0.713 3.766 0.906 ;
      RECT 3.645 0.713 3.656 0.906 ;
      RECT 3.585 0.150 3.645 0.906 ;
      RECT 3.556 0.150 3.585 0.352 ;
      RECT 3.566 0.713 3.585 0.906 ;
      RECT 3.291 0.168 3.556 0.223 ;
      RECT 3.456 0.721 3.467 0.940 ;
      RECT 3.396 0.290 3.456 0.940 ;
      RECT 3.356 0.290 3.396 0.371 ;
      RECT 3.377 0.721 3.396 0.940 ;
      RECT 2.607 0.886 3.377 0.940 ;
      RECT 3.230 0.168 3.291 0.831 ;
      RECT 3.167 0.239 3.230 0.320 ;
      RECT 3.188 0.776 3.230 0.831 ;
      RECT 2.923 0.265 3.167 0.320 ;
      RECT 2.727 0.776 3.066 0.831 ;
      RECT 2.649 0.150 3.018 0.205 ;
      RECT 2.863 0.265 2.923 0.721 ;
      RECT 2.729 0.265 2.863 0.346 ;
      RECT 2.788 0.667 2.863 0.721 ;
      RECT 2.667 0.654 2.727 0.831 ;
      RECT 2.649 0.654 2.667 0.735 ;
      RECT 2.588 0.150 2.649 0.735 ;
      RECT 2.546 0.831 2.607 0.940 ;
      RECT 2.540 0.192 2.588 0.412 ;
      RECT 2.528 0.831 2.546 0.886 ;
      RECT 1.961 0.192 2.540 0.246 ;
      RECT 2.467 0.476 2.528 0.886 ;
      RECT 2.425 0.940 2.486 1.050 ;
      RECT 2.373 0.476 2.467 0.531 ;
      RECT 2.087 0.940 2.425 0.995 ;
      RECT 2.318 0.625 2.407 0.706 ;
      RECT 2.312 0.302 2.373 0.531 ;
      RECT 2.252 0.625 2.318 0.680 ;
      RECT 2.089 0.302 2.312 0.357 ;
      RECT 2.223 0.412 2.252 0.680 ;
      RECT 2.163 0.412 2.223 0.842 ;
      RECT 1.616 0.787 2.163 0.842 ;
      RECT 2.029 0.302 2.089 0.732 ;
      RECT 2.026 0.896 2.087 0.995 ;
      RECT 1.782 0.677 2.029 0.732 ;
      RECT 1.417 0.896 2.026 0.951 ;
      RECT 1.871 0.192 1.961 0.610 ;
      RECT 1.317 0.192 1.871 0.246 ;
      RECT 1.782 0.348 1.811 0.429 ;
      RECT 1.722 0.301 1.782 0.732 ;
      RECT 1.245 0.301 1.722 0.356 ;
      RECT 1.677 0.677 1.722 0.732 ;
      RECT 1.556 0.411 1.616 0.842 ;
      RECT 1.367 0.411 1.556 0.492 ;
      RECT 1.296 0.787 1.556 0.842 ;
      RECT 1.401 0.570 1.430 0.651 ;
      RECT 1.356 0.896 1.417 0.977 ;
      RECT 1.341 0.570 1.401 0.732 ;
      RECT 1.102 0.923 1.356 0.977 ;
      RECT 1.202 0.677 1.341 0.732 ;
      RECT 1.228 0.150 1.317 0.246 ;
      RECT 1.236 0.787 1.296 0.855 ;
      RECT 1.184 0.301 1.245 0.450 ;
      RECT 0.751 0.800 1.236 0.855 ;
      RECT 0.536 0.150 1.228 0.205 ;
      RECT 0.924 0.395 1.184 0.450 ;
      RECT 1.035 0.260 1.124 0.340 ;
      RECT 1.012 0.910 1.102 0.990 ;
      RECT 0.725 0.260 1.035 0.314 ;
      RECT 0.699 0.910 1.012 0.964 ;
      RECT 0.896 0.369 0.924 0.450 ;
      RECT 0.896 0.664 0.902 0.745 ;
      RECT 0.835 0.369 0.896 0.745 ;
      RECT 0.813 0.664 0.835 0.745 ;
      RECT 0.691 0.536 0.751 0.855 ;
      RECT 0.696 0.260 0.725 0.340 ;
      RECT 0.630 0.910 0.699 0.990 ;
      RECT 0.636 0.260 0.696 0.481 ;
      RECT 0.630 0.426 0.636 0.481 ;
      RECT 0.609 0.426 0.630 0.990 ;
      RECT 0.570 0.426 0.609 0.977 ;
      RECT 0.509 0.150 0.536 0.371 ;
      RECT 0.449 0.150 0.509 0.771 ;
      RECT 0.446 0.150 0.449 0.371 ;
      RECT 0.420 0.688 0.449 0.771 ;
      RECT 0.152 0.688 0.420 0.743 ;
      RECT 0.108 0.688 0.152 0.771 ;
      RECT 0.108 0.182 0.137 0.375 ;
      RECT 0.047 0.182 0.108 0.771 ;
  END
END XNOR3X4

MACRO XNOR3X2
  CLASS CORE ;
  FOREIGN XNOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.152 0.227 3.165 0.720 ;
      RECT 3.142 0.199 3.152 0.733 ;
      RECT 3.103 0.199 3.142 0.761 ;
      RECT 3.060 0.199 3.103 0.392 ;
      RECT 3.080 0.652 3.103 0.761 ;
      RECT 3.060 0.652 3.080 0.733 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.672 0.788 2.815 0.900 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.892 0.573 1.898 0.627 ;
      RECT 1.863 0.573 1.892 0.769 ;
      RECT 1.801 0.426 1.863 0.769 ;
      RECT 1.714 0.426 1.801 0.507 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.120 0.526 0.221 0.607 ;
      RECT 0.058 0.526 0.120 0.627 ;
      RECT 0.038 0.526 0.058 0.607 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.947 -0.080 3.200 0.080 ;
      RECT 2.855 -0.080 2.947 0.135 ;
      RECT 0.995 -0.080 2.855 0.080 ;
      RECT 0.904 -0.080 0.995 0.179 ;
      RECT 0.140 -0.080 0.904 0.080 ;
      RECT 0.048 -0.080 0.140 0.359 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.968 1.120 3.200 1.280 ;
      RECT 2.877 0.953 2.968 1.280 ;
      RECT 0.952 1.120 2.877 1.280 ;
      RECT 0.861 1.011 0.952 1.280 ;
      RECT 0.162 1.120 0.861 1.280 ;
      RECT 0.070 0.953 0.162 1.280 ;
      RECT 0.000 1.120 0.070 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.998 0.507 3.041 0.588 ;
      RECT 2.936 0.238 2.998 0.588 ;
      RECT 2.742 0.238 2.936 0.293 ;
      RECT 2.723 0.348 2.785 0.429 ;
      RECT 2.723 0.652 2.774 0.733 ;
      RECT 2.680 0.150 2.742 0.293 ;
      RECT 2.661 0.348 2.723 0.733 ;
      RECT 2.392 0.150 2.680 0.205 ;
      RECT 2.632 0.526 2.661 0.607 ;
      RECT 2.567 0.271 2.597 0.352 ;
      RECT 2.567 0.713 2.586 0.906 ;
      RECT 2.556 0.271 2.567 0.906 ;
      RECT 2.505 0.271 2.556 1.050 ;
      RECT 2.494 0.713 2.505 1.050 ;
      RECT 1.243 0.995 2.494 1.050 ;
      RECT 2.373 0.150 2.392 0.343 ;
      RECT 2.373 0.713 2.392 0.906 ;
      RECT 2.311 0.150 2.373 0.906 ;
      RECT 2.300 0.150 2.311 0.343 ;
      RECT 2.300 0.713 2.311 0.906 ;
      RECT 2.136 0.150 2.198 0.906 ;
      RECT 2.106 0.150 2.136 0.352 ;
      RECT 2.106 0.713 2.136 0.906 ;
      RECT 1.653 0.150 2.106 0.205 ;
      RECT 1.982 0.290 2.044 0.940 ;
      RECT 1.902 0.290 1.982 0.371 ;
      RECT 1.912 0.860 1.982 0.940 ;
      RECT 1.367 0.886 1.912 0.940 ;
      RECT 1.647 0.655 1.739 0.736 ;
      RECT 1.623 0.150 1.653 0.412 ;
      RECT 1.623 0.655 1.647 0.710 ;
      RECT 1.591 0.150 1.623 0.710 ;
      RECT 1.561 0.219 1.591 0.710 ;
      RECT 1.491 0.776 1.545 0.831 ;
      RECT 1.459 0.249 1.491 0.831 ;
      RECT 1.429 0.200 1.459 0.831 ;
      RECT 1.367 0.200 1.429 0.304 ;
      RECT 0.871 0.249 1.367 0.304 ;
      RECT 1.305 0.358 1.367 0.940 ;
      RECT 0.995 0.358 1.305 0.413 ;
      RECT 1.230 0.468 1.243 0.523 ;
      RECT 1.181 0.887 1.243 1.050 ;
      RECT 1.200 0.468 1.230 0.667 ;
      RECT 1.138 0.468 1.200 0.832 ;
      RECT 0.539 0.887 1.181 0.942 ;
      RECT 0.593 0.777 1.138 0.832 ;
      RECT 0.933 0.358 0.995 0.723 ;
      RECT 0.718 0.668 0.933 0.723 ;
      RECT 0.842 0.249 0.871 0.610 ;
      RECT 0.780 0.150 0.842 0.610 ;
      RECT 0.345 0.150 0.780 0.205 ;
      RECT 0.656 0.267 0.718 0.723 ;
      RECT 0.531 0.493 0.593 0.832 ;
      RECT 0.469 0.260 0.539 0.340 ;
      RECT 0.469 0.887 0.539 0.968 ;
      RECT 0.447 0.260 0.469 0.968 ;
      RECT 0.407 0.273 0.447 0.955 ;
      RECT 0.283 0.150 0.345 0.745 ;
      RECT 0.253 0.150 0.283 0.350 ;
      RECT 0.253 0.664 0.283 0.745 ;
  END
END XNOR3X2

MACRO ram_256x16A
  CLASS RING ;
  FOREIGN ram_256x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 59.822 BY 18.924 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.998 1.720 31.108 1.930 ;
      LAYER Metal2 ;
      RECT 30.998 1.720 31.108 1.930 ;
      LAYER Metal3 ;
      RECT 30.998 1.720 31.108 1.930 ;
      LAYER Metal4 ;
      RECT 30.998 1.720 31.108 1.930 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.632 1.720 30.742 1.930 ;
      LAYER Metal2 ;
      RECT 30.632 1.720 30.742 1.930 ;
      LAYER Metal3 ;
      RECT 30.632 1.720 30.742 1.930 ;
      LAYER Metal4 ;
      RECT 30.632 1.720 30.742 1.930 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.118 1.720 30.228 1.930 ;
      LAYER Metal2 ;
      RECT 30.118 1.720 30.228 1.930 ;
      LAYER Metal3 ;
      RECT 30.118 1.720 30.228 1.930 ;
      LAYER Metal4 ;
      RECT 30.118 1.720 30.228 1.930 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 29.752 1.720 29.862 1.930 ;
      LAYER Metal2 ;
      RECT 29.752 1.720 29.862 1.930 ;
      LAYER Metal3 ;
      RECT 29.752 1.720 29.862 1.930 ;
      LAYER Metal4 ;
      RECT 29.752 1.720 29.862 1.930 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 28.872 1.720 28.982 1.930 ;
      LAYER Metal2 ;
      RECT 28.872 1.720 28.982 1.930 ;
      LAYER Metal3 ;
      RECT 28.872 1.720 28.982 1.930 ;
      LAYER Metal4 ;
      RECT 28.872 1.720 28.982 1.930 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 28.358 1.720 28.468 1.930 ;
      LAYER Metal2 ;
      RECT 28.358 1.720 28.468 1.930 ;
      LAYER Metal3 ;
      RECT 28.358 1.720 28.468 1.930 ;
      LAYER Metal4 ;
      RECT 28.358 1.720 28.468 1.930 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.992 1.720 28.102 1.930 ;
      LAYER Metal2 ;
      RECT 27.992 1.720 28.102 1.930 ;
      LAYER Metal3 ;
      RECT 27.992 1.720 28.102 1.930 ;
      LAYER Metal4 ;
      RECT 27.992 1.720 28.102 1.930 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.112 1.720 27.222 1.930 ;
      LAYER Metal2 ;
      RECT 27.112 1.720 27.222 1.930 ;
      LAYER Metal3 ;
      RECT 27.112 1.720 27.222 1.930 ;
      LAYER Metal4 ;
      RECT 27.112 1.720 27.222 1.930 ;
      END
    END A[7]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 31.868 1.720 31.978 1.930 ;
      LAYER Metal2 ;
      RECT 31.868 1.720 31.978 1.930 ;
      LAYER Metal3 ;
      RECT 31.868 1.720 31.978 1.930 ;
      LAYER Metal4 ;
      RECT 31.868 1.720 31.978 1.930 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
      RECT 33.321 1.720 33.431 1.930 ;
      LAYER Metal2 ;
      RECT 33.321 1.720 33.431 1.930 ;
      LAYER Metal3 ;
      RECT 33.321 1.720 33.431 1.930 ;
      LAYER Metal4 ;
      RECT 33.321 1.720 33.431 1.930 ;
      END
    END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal2 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal3 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal4 ;
      RECT 4.546 1.720 4.656 1.930 ;
      END
    END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 41.948 1.720 42.058 1.930 ;
      LAYER Metal2 ;
      RECT 41.948 1.720 42.058 1.930 ;
      LAYER Metal3 ;
      RECT 41.948 1.720 42.058 1.930 ;
      LAYER Metal4 ;
      RECT 41.948 1.720 42.058 1.930 ;
      END
    END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 43.030 1.720 43.140 1.930 ;
      LAYER Metal2 ;
      RECT 43.030 1.720 43.140 1.930 ;
      LAYER Metal3 ;
      RECT 43.030 1.720 43.140 1.930 ;
      LAYER Metal4 ;
      RECT 43.030 1.720 43.140 1.930 ;
      END
    END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 48.016 1.720 48.126 1.930 ;
      LAYER Metal2 ;
      RECT 48.016 1.720 48.126 1.930 ;
      LAYER Metal3 ;
      RECT 48.016 1.720 48.126 1.930 ;
      LAYER Metal4 ;
      RECT 48.016 1.720 48.126 1.930 ;
      END
    END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 49.098 1.720 49.208 1.930 ;
      LAYER Metal2 ;
      RECT 49.098 1.720 49.208 1.930 ;
      LAYER Metal3 ;
      RECT 49.098 1.720 49.208 1.930 ;
      LAYER Metal4 ;
      RECT 49.098 1.720 49.208 1.930 ;
      END
    END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 54.084 1.720 54.194 1.930 ;
      LAYER Metal2 ;
      RECT 54.084 1.720 54.194 1.930 ;
      LAYER Metal3 ;
      RECT 54.084 1.720 54.194 1.930 ;
      LAYER Metal4 ;
      RECT 54.084 1.720 54.194 1.930 ;
      END
    END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 55.166 1.720 55.276 1.930 ;
      LAYER Metal2 ;
      RECT 55.166 1.720 55.276 1.930 ;
      LAYER Metal3 ;
      RECT 55.166 1.720 55.276 1.930 ;
      LAYER Metal4 ;
      RECT 55.166 1.720 55.276 1.930 ;
      END
    END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal2 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal3 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal4 ;
      RECT 5.628 1.720 5.738 1.930 ;
      END
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal2 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal3 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal4 ;
      RECT 10.614 1.720 10.724 1.930 ;
      END
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal2 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal3 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal4 ;
      RECT 11.696 1.720 11.806 1.930 ;
      END
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal2 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal3 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal4 ;
      RECT 16.682 1.720 16.792 1.930 ;
      END
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal2 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal3 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal4 ;
      RECT 17.764 1.720 17.874 1.930 ;
      END
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal2 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal3 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal4 ;
      RECT 22.750 1.720 22.860 1.930 ;
      END
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal2 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal3 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal4 ;
      RECT 23.832 1.720 23.942 1.930 ;
      END
    END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 35.880 1.720 35.990 1.930 ;
      LAYER Metal2 ;
      RECT 35.880 1.720 35.990 1.930 ;
      LAYER Metal3 ;
      RECT 35.880 1.720 35.990 1.930 ;
      LAYER Metal4 ;
      RECT 35.880 1.720 35.990 1.930 ;
      END
    END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 36.962 1.720 37.072 1.930 ;
      LAYER Metal2 ;
      RECT 36.962 1.720 37.072 1.930 ;
      LAYER Metal3 ;
      RECT 36.962 1.720 37.072 1.930 ;
      LAYER Metal4 ;
      RECT 36.962 1.720 37.072 1.930 ;
      END
    END D[9]
  PIN OEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 33.020 1.720 33.130 1.930 ;
      LAYER Metal2 ;
      RECT 33.020 1.720 33.130 1.930 ;
      LAYER Metal3 ;
      RECT 33.020 1.720 33.130 1.930 ;
      LAYER Metal4 ;
      RECT 33.020 1.720 33.130 1.930 ;
      END
    END OEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal2 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal3 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal4 ;
      RECT 3.998 1.720 4.108 1.930 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 41.420 1.720 41.530 1.930 ;
      LAYER Metal2 ;
      RECT 41.420 1.720 41.530 1.930 ;
      LAYER Metal3 ;
      RECT 41.420 1.720 41.530 1.930 ;
      LAYER Metal4 ;
      RECT 41.420 1.720 41.530 1.930 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 43.558 1.720 43.668 1.930 ;
      LAYER Metal2 ;
      RECT 43.558 1.720 43.668 1.930 ;
      LAYER Metal3 ;
      RECT 43.558 1.720 43.668 1.930 ;
      LAYER Metal4 ;
      RECT 43.558 1.720 43.668 1.930 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 47.488 1.720 47.598 1.930 ;
      LAYER Metal2 ;
      RECT 47.488 1.720 47.598 1.930 ;
      LAYER Metal3 ;
      RECT 47.488 1.720 47.598 1.930 ;
      LAYER Metal4 ;
      RECT 47.488 1.720 47.598 1.930 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 49.626 1.720 49.736 1.930 ;
      LAYER Metal2 ;
      RECT 49.626 1.720 49.736 1.930 ;
      LAYER Metal3 ;
      RECT 49.626 1.720 49.736 1.930 ;
      LAYER Metal4 ;
      RECT 49.626 1.720 49.736 1.930 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 53.556 1.720 53.666 1.930 ;
      LAYER Metal2 ;
      RECT 53.556 1.720 53.666 1.930 ;
      LAYER Metal3 ;
      RECT 53.556 1.720 53.666 1.930 ;
      LAYER Metal4 ;
      RECT 53.556 1.720 53.666 1.930 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 55.704 1.720 55.814 1.930 ;
      LAYER Metal2 ;
      RECT 55.704 1.720 55.814 1.930 ;
      LAYER Metal3 ;
      RECT 55.704 1.720 55.814 1.930 ;
      LAYER Metal4 ;
      RECT 55.704 1.720 55.814 1.930 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal2 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal3 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal4 ;
      RECT 6.156 1.720 6.266 1.930 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal2 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal3 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal4 ;
      RECT 10.086 1.720 10.196 1.930 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal2 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal3 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal4 ;
      RECT 12.224 1.720 12.334 1.930 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal2 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal3 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal4 ;
      RECT 16.154 1.720 16.264 1.930 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal2 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal3 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal4 ;
      RECT 18.292 1.720 18.402 1.930 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal2 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal3 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal4 ;
      RECT 22.222 1.720 22.332 1.930 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal2 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal3 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal4 ;
      RECT 24.360 1.720 24.470 1.930 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 35.352 1.720 35.462 1.930 ;
      LAYER Metal2 ;
      RECT 35.352 1.720 35.462 1.930 ;
      LAYER Metal3 ;
      RECT 35.352 1.720 35.462 1.930 ;
      LAYER Metal4 ;
      RECT 35.352 1.720 35.462 1.930 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 37.490 1.720 37.600 1.930 ;
      LAYER Metal2 ;
      RECT 37.490 1.720 37.600 1.930 ;
      LAYER Metal3 ;
      RECT 37.490 1.720 37.600 1.930 ;
      LAYER Metal4 ;
      RECT 37.490 1.720 37.600 1.930 ;
      END
    END Q[9]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 32.156 1.720 32.266 1.930 ;
      LAYER Metal2 ;
      RECT 32.156 1.720 32.266 1.930 ;
      LAYER Metal3 ;
      RECT 32.156 1.720 32.266 1.930 ;
      LAYER Metal4 ;
      RECT 32.156 1.720 32.266 1.930 ;
      END
    END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.000 18.224 59.822 18.924 ;
      LAYER Metal5 ;
      RECT 0.000 0.000 59.822 0.700 ;
      LAYER Metal4 ;
      RECT 59.122 0.000 59.822 18.924 ;
      LAYER Metal4 ;
      RECT 0.000 0.000 0.700 18.924 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.860 17.364 58.962 18.064 ;
      LAYER Metal5 ;
      RECT 0.860 0.860 58.962 1.560 ;
      LAYER Metal4 ;
      RECT 58.262 0.860 58.962 18.064 ;
      LAYER Metal4 ;
      RECT 0.860 0.860 1.560 18.064 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 1.720 1.720 58.102 17.204 ;
    LAYER Metal1 ;
    RECT 1.720 1.980 58.102 17.204 ;
    RECT 1.720 1.720 3.898 17.204 ;
    RECT 55.840 1.720 58.102 17.204 ;
    LAYER Metal2 ;
    RECT 1.720 1.980 58.102 17.204 ;
    RECT 1.720 1.720 3.898 17.204 ;
    RECT 55.840 1.720 58.102 17.204 ;
    LAYER Metal3 ;
    RECT 1.720 1.980 58.102 17.204 ;
    RECT 1.720 1.720 3.898 17.204 ;
    RECT 55.840 1.720 58.102 17.204 ;
    LAYER Metal4 ;
    RECT 1.720 1.980 58.102 17.204 ;
    RECT 1.720 1.720 3.898 17.204 ;
    RECT 55.840 1.720 58.102 17.204 ;
    LAYER Via1 ;
    RECT 1.720 1.720 58.102 17.204 ;
    LAYER Via2 ;
    RECT 1.720 1.720 58.102 17.204 ;
    LAYER Via3 ;
    RECT 1.720 1.720 58.102 17.204 ;
    END
END ram_256x16A

MACRO rom_512x16A
  CLASS RING ;
  FOREIGN rom_512x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 36.817 BY 18.684 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 8.870 2.120 8.981 2.330 ;
      LAYER Metal2 ;
      RECT 8.870 2.120 8.981 2.330 ;
      LAYER Metal3 ;
      RECT 8.870 2.120 8.981 2.330 ;
      LAYER Metal4 ;
      RECT 8.870 2.120 8.981 2.330 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 8.421 2.120 8.531 2.330 ;
      LAYER Metal2 ;
      RECT 8.421 2.120 8.531 2.330 ;
      LAYER Metal3 ;
      RECT 8.421 2.120 8.531 2.330 ;
      LAYER Metal4 ;
      RECT 8.421 2.120 8.531 2.330 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 7.971 2.120 8.081 2.330 ;
      LAYER Metal2 ;
      RECT 7.971 2.120 8.081 2.330 ;
      LAYER Metal3 ;
      RECT 7.971 2.120 8.081 2.330 ;
      LAYER Metal4 ;
      RECT 7.971 2.120 8.081 2.330 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 7.071 2.120 7.181 2.330 ;
      LAYER Metal2 ;
      RECT 7.071 2.120 7.181 2.330 ;
      LAYER Metal3 ;
      RECT 7.071 2.120 7.181 2.330 ;
      LAYER Metal4 ;
      RECT 7.071 2.120 7.181 2.330 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 6.171 2.120 6.281 2.330 ;
      LAYER Metal2 ;
      RECT 6.171 2.120 6.281 2.330 ;
      LAYER Metal3 ;
      RECT 6.171 2.120 6.281 2.330 ;
      LAYER Metal4 ;
      RECT 6.171 2.120 6.281 2.330 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 5.721 2.120 5.831 2.330 ;
      LAYER Metal2 ;
      RECT 5.721 2.120 5.831 2.330 ;
      LAYER Metal3 ;
      RECT 5.721 2.120 5.831 2.330 ;
      LAYER Metal4 ;
      RECT 5.721 2.120 5.831 2.330 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 5.271 2.120 5.381 2.330 ;
      LAYER Metal2 ;
      RECT 5.271 2.120 5.381 2.330 ;
      LAYER Metal3 ;
      RECT 5.271 2.120 5.381 2.330 ;
      LAYER Metal4 ;
      RECT 5.271 2.120 5.381 2.330 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 4.370 2.120 4.481 2.330 ;
      LAYER Metal2 ;
      RECT 4.370 2.120 4.481 2.330 ;
      LAYER Metal3 ;
      RECT 4.370 2.120 4.481 2.330 ;
      LAYER Metal4 ;
      RECT 4.370 2.120 4.481 2.330 ;
      END
    END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 3.921 2.120 4.030 2.330 ;
      LAYER Metal2 ;
      RECT 3.921 2.120 4.030 2.330 ;
      LAYER Metal3 ;
      RECT 3.921 2.120 4.030 2.330 ;
      LAYER Metal4 ;
      RECT 3.921 2.120 4.030 2.330 ;
      END
    END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 11.202 2.120 11.312 2.330 ;
      LAYER Metal2 ;
      RECT 11.202 2.120 11.312 2.330 ;
      LAYER Metal3 ;
      RECT 11.202 2.120 11.312 2.330 ;
      LAYER Metal4 ;
      RECT 11.202 2.120 11.312 2.330 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
      RECT 11.032 2.120 11.142 2.330 ;
      LAYER Metal2 ;
      RECT 11.032 2.120 11.142 2.330 ;
      LAYER Metal3 ;
      RECT 11.032 2.120 11.142 2.330 ;
      LAYER Metal4 ;
      RECT 11.032 2.120 11.142 2.330 ;
      END
    END CLK
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 14.157 2.120 14.268 2.330 ;
      LAYER Metal2 ;
      RECT 14.157 2.120 14.268 2.330 ;
      LAYER Metal3 ;
      RECT 14.157 2.120 14.268 2.330 ;
      LAYER Metal4 ;
      RECT 14.157 2.120 14.268 2.330 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.548 2.120 27.657 2.330 ;
      LAYER Metal2 ;
      RECT 27.548 2.120 27.657 2.330 ;
      LAYER Metal3 ;
      RECT 27.548 2.120 27.657 2.330 ;
      LAYER Metal4 ;
      RECT 27.548 2.120 27.657 2.330 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.854 2.120 27.963 2.330 ;
      LAYER Metal2 ;
      RECT 27.854 2.120 27.963 2.330 ;
      LAYER Metal3 ;
      RECT 27.854 2.120 27.963 2.330 ;
      LAYER Metal4 ;
      RECT 27.854 2.120 27.963 2.330 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.226 2.120 30.336 2.330 ;
      LAYER Metal2 ;
      RECT 30.226 2.120 30.336 2.330 ;
      LAYER Metal3 ;
      RECT 30.226 2.120 30.336 2.330 ;
      LAYER Metal4 ;
      RECT 30.226 2.120 30.336 2.330 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.532 2.120 30.642 2.330 ;
      LAYER Metal2 ;
      RECT 30.532 2.120 30.642 2.330 ;
      LAYER Metal3 ;
      RECT 30.532 2.120 30.642 2.330 ;
      LAYER Metal4 ;
      RECT 30.532 2.120 30.642 2.330 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 32.904 2.120 33.014 2.330 ;
      LAYER Metal2 ;
      RECT 32.904 2.120 33.014 2.330 ;
      LAYER Metal3 ;
      RECT 32.904 2.120 33.014 2.330 ;
      LAYER Metal4 ;
      RECT 32.904 2.120 33.014 2.330 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 33.210 2.120 33.320 2.330 ;
      LAYER Metal2 ;
      RECT 33.210 2.120 33.320 2.330 ;
      LAYER Metal3 ;
      RECT 33.210 2.120 33.320 2.330 ;
      LAYER Metal4 ;
      RECT 33.210 2.120 33.320 2.330 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 14.463 2.120 14.574 2.330 ;
      LAYER Metal2 ;
      RECT 14.463 2.120 14.574 2.330 ;
      LAYER Metal3 ;
      RECT 14.463 2.120 14.574 2.330 ;
      LAYER Metal4 ;
      RECT 14.463 2.120 14.574 2.330 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 16.835 2.120 16.946 2.330 ;
      LAYER Metal2 ;
      RECT 16.835 2.120 16.946 2.330 ;
      LAYER Metal3 ;
      RECT 16.835 2.120 16.946 2.330 ;
      LAYER Metal4 ;
      RECT 16.835 2.120 16.946 2.330 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 17.142 2.120 17.252 2.330 ;
      LAYER Metal2 ;
      RECT 17.142 2.120 17.252 2.330 ;
      LAYER Metal3 ;
      RECT 17.142 2.120 17.252 2.330 ;
      LAYER Metal4 ;
      RECT 17.142 2.120 17.252 2.330 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 19.514 2.120 19.624 2.330 ;
      LAYER Metal2 ;
      RECT 19.514 2.120 19.624 2.330 ;
      LAYER Metal3 ;
      RECT 19.514 2.120 19.624 2.330 ;
      LAYER Metal4 ;
      RECT 19.514 2.120 19.624 2.330 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 19.820 2.120 19.930 2.330 ;
      LAYER Metal2 ;
      RECT 19.820 2.120 19.930 2.330 ;
      LAYER Metal3 ;
      RECT 19.820 2.120 19.930 2.330 ;
      LAYER Metal4 ;
      RECT 19.820 2.120 19.930 2.330 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.192 2.120 22.302 2.330 ;
      LAYER Metal2 ;
      RECT 22.192 2.120 22.302 2.330 ;
      LAYER Metal3 ;
      RECT 22.192 2.120 22.302 2.330 ;
      LAYER Metal4 ;
      RECT 22.192 2.120 22.302 2.330 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.498 2.120 22.608 2.330 ;
      LAYER Metal2 ;
      RECT 22.498 2.120 22.608 2.330 ;
      LAYER Metal3 ;
      RECT 22.498 2.120 22.608 2.330 ;
      LAYER Metal4 ;
      RECT 22.498 2.120 22.608 2.330 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 24.870 2.120 24.980 2.330 ;
      LAYER Metal2 ;
      RECT 24.870 2.120 24.980 2.330 ;
      LAYER Metal3 ;
      RECT 24.870 2.120 24.980 2.330 ;
      LAYER Metal4 ;
      RECT 24.870 2.120 24.980 2.330 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 25.175 2.120 25.285 2.330 ;
      LAYER Metal2 ;
      RECT 25.175 2.120 25.285 2.330 ;
      LAYER Metal3 ;
      RECT 25.175 2.120 25.285 2.330 ;
      LAYER Metal4 ;
      RECT 25.175 2.120 25.285 2.330 ;
      END
    END Q[9]
  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.000 17.784 36.817 18.684 ;
      LAYER Metal5 ;
      RECT 0.000 0.000 36.817 0.900 ;
      LAYER Metal4 ;
      RECT 35.917 0.000 36.817 18.684 ;
      LAYER Metal4 ;
      RECT 0.000 0.000 0.900 18.684 ;
      END
    END VDD
  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 1.060 16.725 35.757 17.625 ;
      LAYER Metal5 ;
      RECT 1.060 1.060 35.757 1.960 ;
      LAYER Metal4 ;
      RECT 34.857 1.060 35.757 17.625 ;
      LAYER Metal4 ;
      RECT 1.060 1.060 1.960 17.625 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 2.120 2.120 34.697 16.565 ;
    LAYER Metal1 ;
    RECT 2.120 2.380 34.697 16.565 ;
    RECT 2.120 2.120 3.821 16.565 ;
    RECT 33.310 2.380 34.697 16.565 ;
    LAYER Metal2 ;
    RECT 2.120 2.380 34.697 16.565 ;
    RECT 2.120 2.120 3.821 16.565 ;
    RECT 33.310 2.380 34.697 16.565 ;
    LAYER Metal3 ;
    RECT 2.120 2.380 34.697 16.565 ;
    RECT 2.120 2.120 3.821 16.565 ;
    RECT 33.310 2.380 34.697 16.565 ;
    LAYER Metal4 ;
    RECT 2.120 2.380 34.697 16.565 ;
    RECT 2.120 2.120 3.821 16.565 ;
    RECT 33.310 2.380 34.697 16.565 ;
    LAYER Via1 ;
    RECT 2.120 2.120 34.697 16.565 ;
    LAYER Via2 ;
    RECT 2.120 2.120 34.697 16.565 ;
    LAYER Via3 ;
    RECT 2.120 2.120 34.697 16.565 ;
    END
END rom_512x16A

MACRO pllclk
  CLASS BLOCK ;
  ORIGIN 0.06 0 ;
  SIZE 15.006 BY 27.359 ;
  SYMMETRY X Y R90 ;

  PIN refclk
  DIRECTION INPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 15.000 0.260 15.200 ;
      LAYER Metal3 ;
      RECT 0.000 15.000 0.260 15.200 ;
     END
  END refclk

  PIN clk1x
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 5.000 0.260 5.200 ;
      LAYER Metal3 ;
      RECT 0.000 5.000 0.260 5.200 ;
     END
  END clk1x

  PIN clk2x
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 6.000 0.260 6.200 ;
      LAYER Metal3 ;
      RECT 0.000 6.000 0.260 6.200 ;
     END
  END clk2x

  PIN ibias
  DIRECTION INPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 18.040 0.260 18.190 ;
      LAYER Metal3 ;
      RECT 0.000 18.040 0.260 18.190 ;
     END
  END ibias

  PIN reset
  DIRECTION INPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 18.504 0.260 18.654 ;
      LAYER Metal3 ;
      RECT 0.000 18.504 0.260 18.654 ;
     END
  END reset

  PIN vcom
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 17.122 0.260 17.272 ;
      LAYER Metal3 ;
      RECT 0.000 17.122 0.260 17.272 ;
     END
  END vcom

  PIN vcop
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal2 ;
      RECT 0.000 17.586 0.260 17.736 ;
      LAYER Metal3 ;
      RECT 0.000 17.586 0.260 17.736 ;
     END
  END vcop

  PIN AVSS
  DIRECTION INOUT ;
  USE GROUND ;
     PORT
      LAYER Metal3 ;
      RECT 14.740 17.846 15.000 18.346 ;
     END
  END AVSS

  PIN AVDD
  DIRECTION INOUT ;
  USE POWER ;
     PORT
      LAYER Metal3 ;
      RECT 14.740 16.185 15.000 16.686 ;
     END
  END AVDD
  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
     PORT
      LAYER Metal3 ;
      RECT 14.740 2.137 15.000 2.637 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
     PORT
      LAYER Metal3 ;
      RECT 14.740 0.477 15.000 0.977 ;
     END
  END VDD
  OBS
      LAYER OVERLAP ;
	RECT 0.000 0.000 15.006 27.359 ;
      LAYER Metal1 ;
	RECT 0.000 0.000 15.006 27.359 ;
      LAYER Metal2 ;
	RECT 0.310 0.000 15.006 27.359 ;
	RECT 0.000 0.000 15.006 4.500 ;
	RECT 0.000 19.100 15.006 27.359 ;
	RECT 0.000 6.700 15.006 14.500 ;
      LAYER Metal3 ;
	RECT 0.310 0.000 14.690 27.359 ;
	RECT 0.000 0.000 14.690 4.500 ;
	RECT 0.000 19.100 14.690 27.359 ;
	RECT 0.000 6.700 14.690 14.500 ;
      LAYER Metal4 ;
	RECT 0.000 0.000 15.006 27.359 ;
      LAYER Metal5 ;
	RECT 0.000 0.000 15.006 27.359 ;
      LAYER Metal6 ;
	RECT 0.000 0.000 15.006 27.359 ;
  END
END pllclk

MACRO ram_128x16A
  CLASS RING ;
  FOREIGN ram_128x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 59.382 BY 16.899 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.558 1.720 30.668 1.930 ;
      LAYER Metal2 ;
      RECT 30.558 1.720 30.668 1.930 ;
      LAYER Metal3 ;
      RECT 30.558 1.720 30.668 1.930 ;
      LAYER Metal4 ;
      RECT 30.558 1.720 30.668 1.930 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 30.192 1.720 30.302 1.930 ;
      LAYER Metal2 ;
      RECT 30.192 1.720 30.302 1.930 ;
      LAYER Metal3 ;
      RECT 30.192 1.720 30.302 1.930 ;
      LAYER Metal4 ;
      RECT 30.192 1.720 30.302 1.930 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 29.678 1.720 29.788 1.930 ;
      LAYER Metal2 ;
      RECT 29.678 1.720 29.788 1.930 ;
      LAYER Metal3 ;
      RECT 29.678 1.720 29.788 1.930 ;
      LAYER Metal4 ;
      RECT 29.678 1.720 29.788 1.930 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 29.312 1.720 29.422 1.930 ;
      LAYER Metal2 ;
      RECT 29.312 1.720 29.422 1.930 ;
      LAYER Metal3 ;
      RECT 29.312 1.720 29.422 1.930 ;
      LAYER Metal4 ;
      RECT 29.312 1.720 29.422 1.930 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 28.432 1.720 28.542 1.930 ;
      LAYER Metal2 ;
      RECT 28.432 1.720 28.542 1.930 ;
      LAYER Metal3 ;
      RECT 28.432 1.720 28.542 1.930 ;
      LAYER Metal4 ;
      RECT 28.432 1.720 28.542 1.930 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.918 1.720 28.028 1.930 ;
      LAYER Metal2 ;
      RECT 27.918 1.720 28.028 1.930 ;
      LAYER Metal3 ;
      RECT 27.918 1.720 28.028 1.930 ;
      LAYER Metal4 ;
      RECT 27.918 1.720 28.028 1.930 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 27.552 1.720 27.662 1.930 ;
      LAYER Metal2 ;
      RECT 27.552 1.720 27.662 1.930 ;
      LAYER Metal3 ;
      RECT 27.552 1.720 27.662 1.930 ;
      LAYER Metal4 ;
      RECT 27.552 1.720 27.662 1.930 ;
      END
    END A[6]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 31.428 1.720 31.538 1.930 ;
      LAYER Metal2 ;
      RECT 31.428 1.720 31.538 1.930 ;
      LAYER Metal3 ;
      RECT 31.428 1.720 31.538 1.930 ;
      LAYER Metal4 ;
      RECT 31.428 1.720 31.538 1.930 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
      RECT 32.881 1.720 32.991 1.930 ;
      LAYER Metal2 ;
      RECT 32.881 1.720 32.991 1.930 ;
      LAYER Metal3 ;
      RECT 32.881 1.720 32.991 1.930 ;
      LAYER Metal4 ;
      RECT 32.881 1.720 32.991 1.930 ;
      END
    END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal2 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal3 ;
      RECT 4.546 1.720 4.656 1.930 ;
      LAYER Metal4 ;
      RECT 4.546 1.720 4.656 1.930 ;
      END
    END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 41.508 1.720 41.618 1.930 ;
      LAYER Metal2 ;
      RECT 41.508 1.720 41.618 1.930 ;
      LAYER Metal3 ;
      RECT 41.508 1.720 41.618 1.930 ;
      LAYER Metal4 ;
      RECT 41.508 1.720 41.618 1.930 ;
      END
    END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 42.590 1.720 42.700 1.930 ;
      LAYER Metal2 ;
      RECT 42.590 1.720 42.700 1.930 ;
      LAYER Metal3 ;
      RECT 42.590 1.720 42.700 1.930 ;
      LAYER Metal4 ;
      RECT 42.590 1.720 42.700 1.930 ;
      END
    END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 47.576 1.720 47.686 1.930 ;
      LAYER Metal2 ;
      RECT 47.576 1.720 47.686 1.930 ;
      LAYER Metal3 ;
      RECT 47.576 1.720 47.686 1.930 ;
      LAYER Metal4 ;
      RECT 47.576 1.720 47.686 1.930 ;
      END
    END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 48.658 1.720 48.768 1.930 ;
      LAYER Metal2 ;
      RECT 48.658 1.720 48.768 1.930 ;
      LAYER Metal3 ;
      RECT 48.658 1.720 48.768 1.930 ;
      LAYER Metal4 ;
      RECT 48.658 1.720 48.768 1.930 ;
      END
    END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 53.644 1.720 53.754 1.930 ;
      LAYER Metal2 ;
      RECT 53.644 1.720 53.754 1.930 ;
      LAYER Metal3 ;
      RECT 53.644 1.720 53.754 1.930 ;
      LAYER Metal4 ;
      RECT 53.644 1.720 53.754 1.930 ;
      END
    END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 54.726 1.720 54.836 1.930 ;
      LAYER Metal2 ;
      RECT 54.726 1.720 54.836 1.930 ;
      LAYER Metal3 ;
      RECT 54.726 1.720 54.836 1.930 ;
      LAYER Metal4 ;
      RECT 54.726 1.720 54.836 1.930 ;
      END
    END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal2 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal3 ;
      RECT 5.628 1.720 5.738 1.930 ;
      LAYER Metal4 ;
      RECT 5.628 1.720 5.738 1.930 ;
      END
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal2 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal3 ;
      RECT 10.614 1.720 10.724 1.930 ;
      LAYER Metal4 ;
      RECT 10.614 1.720 10.724 1.930 ;
      END
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal2 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal3 ;
      RECT 11.696 1.720 11.806 1.930 ;
      LAYER Metal4 ;
      RECT 11.696 1.720 11.806 1.930 ;
      END
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal2 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal3 ;
      RECT 16.682 1.720 16.792 1.930 ;
      LAYER Metal4 ;
      RECT 16.682 1.720 16.792 1.930 ;
      END
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal2 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal3 ;
      RECT 17.764 1.720 17.874 1.930 ;
      LAYER Metal4 ;
      RECT 17.764 1.720 17.874 1.930 ;
      END
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal2 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal3 ;
      RECT 22.750 1.720 22.860 1.930 ;
      LAYER Metal4 ;
      RECT 22.750 1.720 22.860 1.930 ;
      END
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal2 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal3 ;
      RECT 23.832 1.720 23.942 1.930 ;
      LAYER Metal4 ;
      RECT 23.832 1.720 23.942 1.930 ;
      END
    END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 35.440 1.720 35.550 1.930 ;
      LAYER Metal2 ;
      RECT 35.440 1.720 35.550 1.930 ;
      LAYER Metal3 ;
      RECT 35.440 1.720 35.550 1.930 ;
      LAYER Metal4 ;
      RECT 35.440 1.720 35.550 1.930 ;
      END
    END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 36.522 1.720 36.632 1.930 ;
      LAYER Metal2 ;
      RECT 36.522 1.720 36.632 1.930 ;
      LAYER Metal3 ;
      RECT 36.522 1.720 36.632 1.930 ;
      LAYER Metal4 ;
      RECT 36.522 1.720 36.632 1.930 ;
      END
    END D[9]
  PIN OEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 32.580 1.720 32.690 1.930 ;
      LAYER Metal2 ;
      RECT 32.580 1.720 32.690 1.930 ;
      LAYER Metal3 ;
      RECT 32.580 1.720 32.690 1.930 ;
      LAYER Metal4 ;
      RECT 32.580 1.720 32.690 1.930 ;
      END
    END OEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal2 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal3 ;
      RECT 3.998 1.720 4.108 1.930 ;
      LAYER Metal4 ;
      RECT 3.998 1.720 4.108 1.930 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 40.980 1.720 41.090 1.930 ;
      LAYER Metal2 ;
      RECT 40.980 1.720 41.090 1.930 ;
      LAYER Metal3 ;
      RECT 40.980 1.720 41.090 1.930 ;
      LAYER Metal4 ;
      RECT 40.980 1.720 41.090 1.930 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 43.118 1.720 43.228 1.930 ;
      LAYER Metal2 ;
      RECT 43.118 1.720 43.228 1.930 ;
      LAYER Metal3 ;
      RECT 43.118 1.720 43.228 1.930 ;
      LAYER Metal4 ;
      RECT 43.118 1.720 43.228 1.930 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 47.048 1.720 47.158 1.930 ;
      LAYER Metal2 ;
      RECT 47.048 1.720 47.158 1.930 ;
      LAYER Metal3 ;
      RECT 47.048 1.720 47.158 1.930 ;
      LAYER Metal4 ;
      RECT 47.048 1.720 47.158 1.930 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 49.186 1.720 49.296 1.930 ;
      LAYER Metal2 ;
      RECT 49.186 1.720 49.296 1.930 ;
      LAYER Metal3 ;
      RECT 49.186 1.720 49.296 1.930 ;
      LAYER Metal4 ;
      RECT 49.186 1.720 49.296 1.930 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 53.116 1.720 53.226 1.930 ;
      LAYER Metal2 ;
      RECT 53.116 1.720 53.226 1.930 ;
      LAYER Metal3 ;
      RECT 53.116 1.720 53.226 1.930 ;
      LAYER Metal4 ;
      RECT 53.116 1.720 53.226 1.930 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 55.264 1.720 55.374 1.930 ;
      LAYER Metal2 ;
      RECT 55.264 1.720 55.374 1.930 ;
      LAYER Metal3 ;
      RECT 55.264 1.720 55.374 1.930 ;
      LAYER Metal4 ;
      RECT 55.264 1.720 55.374 1.930 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal2 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal3 ;
      RECT 6.156 1.720 6.266 1.930 ;
      LAYER Metal4 ;
      RECT 6.156 1.720 6.266 1.930 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal2 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal3 ;
      RECT 10.086 1.720 10.196 1.930 ;
      LAYER Metal4 ;
      RECT 10.086 1.720 10.196 1.930 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal2 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal3 ;
      RECT 12.224 1.720 12.334 1.930 ;
      LAYER Metal4 ;
      RECT 12.224 1.720 12.334 1.930 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal2 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal3 ;
      RECT 16.154 1.720 16.264 1.930 ;
      LAYER Metal4 ;
      RECT 16.154 1.720 16.264 1.930 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal2 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal3 ;
      RECT 18.292 1.720 18.402 1.930 ;
      LAYER Metal4 ;
      RECT 18.292 1.720 18.402 1.930 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal2 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal3 ;
      RECT 22.222 1.720 22.332 1.930 ;
      LAYER Metal4 ;
      RECT 22.222 1.720 22.332 1.930 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal2 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal3 ;
      RECT 24.360 1.720 24.470 1.930 ;
      LAYER Metal4 ;
      RECT 24.360 1.720 24.470 1.930 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 34.912 1.720 35.022 1.930 ;
      LAYER Metal2 ;
      RECT 34.912 1.720 35.022 1.930 ;
      LAYER Metal3 ;
      RECT 34.912 1.720 35.022 1.930 ;
      LAYER Metal4 ;
      RECT 34.912 1.720 35.022 1.930 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 37.050 1.720 37.160 1.930 ;
      LAYER Metal2 ;
      RECT 37.050 1.720 37.160 1.930 ;
      LAYER Metal3 ;
      RECT 37.050 1.720 37.160 1.930 ;
      LAYER Metal4 ;
      RECT 37.050 1.720 37.160 1.930 ;
      END
    END Q[9]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 31.716 1.720 31.826 1.930 ;
      LAYER Metal2 ;
      RECT 31.716 1.720 31.826 1.930 ;
      LAYER Metal3 ;
      RECT 31.716 1.720 31.826 1.930 ;
      LAYER Metal4 ;
      RECT 31.716 1.720 31.826 1.930 ;
      END
    END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.000 16.200 59.382 16.900 ;
      LAYER Metal5 ;
      RECT 0.000 0.000 59.382 0.700 ;
      LAYER Metal4 ;
      RECT 58.682 0.000 59.382 16.899 ;
      LAYER Metal4 ;
      RECT 0.000 0.000 0.700 16.899 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.860 15.340 58.522 16.040 ;
      LAYER Metal5 ;
      RECT 0.860 0.860 58.522 1.560 ;
      LAYER Metal4 ;
      RECT 57.822 0.860 58.522 16.040 ;
      LAYER Metal4 ;
      RECT 0.860 0.860 1.560 16.040 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 1.720 1.720 57.662 15.180 ;
    LAYER Metal1 ;
    RECT 1.720 1.980 57.662 15.180 ;
    RECT 1.720 1.720 3.898 15.180 ;
    RECT 55.474 1.720 57.662 15.180 ;
    LAYER Metal2 ;
    RECT 1.720 1.980 57.662 15.180 ;
    RECT 1.720 1.720 3.898 15.180 ;
    RECT 55.474 1.720 57.662 15.180 ;
    LAYER Metal3 ;
    RECT 1.720 1.980 57.662 15.180 ;
    RECT 1.720 1.720 3.898 15.180 ;
    RECT 55.474 1.720 57.662 15.180 ;
    LAYER Metal4 ;
    RECT 1.720 1.980 57.662 15.180 ;
    RECT 1.720 1.720 3.898 15.180 ;
    RECT 55.474 1.720 57.662 15.180 ;
    LAYER Via1 ;
    RECT 1.720 1.720 57.662 15.180 ;
    LAYER Via2 ;
    RECT 1.720 1.720 57.662 15.180 ;
    LAYER Via3 ;
    RECT 1.720 1.720 57.662 15.180 ;
    END
END ram_128x16A

MACRO PCORNERDG
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNERDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.500 BY 23.500 ;
    SYMMETRY x y r90 ;
    SITE CoreSite ;
    OBS
        LAYER Metal1 ;
        RECT 0.000 0.000 23.500 23.500 ;
        LAYER Metal2 ;
        RECT 0.000 0.000 23.500 23.500 ;
        LAYER Metal3 ;
        RECT 0.000 0.000 23.500 23.500 ;
        LAYER Metal4 ;
        RECT 0.000 0.000 23.500 23.500 ;
        LAYER Metal5 ;
        RECT 0.000 0.000 23.500 23.500 ;
        LAYER Metal6 ;
        RECT 0.000 0.000 23.500 23.500 ;
    END
END PCORNERDG

MACRO PDIDGZ
    CLASS PAD ;
    FOREIGN PDIDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 23.500 ;
    SYMMETRY x y r90 ;
    SITE CoreSite ;
    PIN PAD
        DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT 1.877 0.000 2.224 0.136 ;
        LAYER Metal2 ;
        RECT 1.877 0.000 2.224 0.136 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal2 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal3 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal4 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal5 ;
        RECT 3.217 23.400 3.417 23.500 ;
        END
    END C
    OBS
        LAYER Metal1 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 2.274 0.000 3.167 23.500 ;
        RECT 1.827 0.196 2.274 23.500 ;
        RECT 0.000 0.000 1.827 23.500 ;
        LAYER Via1 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal2 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 2.274 0.000 3.167 23.500 ;
        RECT 1.827 0.196 2.274 23.500 ;
        RECT 0.000 0.000 1.827 23.500 ;
        LAYER Via2 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal3 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via3 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal4 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via4 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal5 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via5 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal6 ;
        RECT 0.000 0.000 4.000 23.500 ;
    END
END PDIDGZ

MACRO PDO04CDG
    CLASS PAD ;
    FOREIGN PDO04CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 23.500 ;
    SYMMETRY x y r90 ;
    SITE CoreSite ;
    PIN PAD
        DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT 1.877 0.000 2.224 0.136 ;
        LAYER Metal2 ;
        RECT 1.877 0.000 2.224 0.136 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal2 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal3 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal4 ;
        RECT 3.217 23.400 3.417 23.500 ;
        LAYER Metal5 ;
        RECT 3.217 23.400 3.417 23.500 ;
        END
    END I
    OBS
        LAYER Metal1 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 2.274 0.000 3.167 23.500 ;
        RECT 1.827 0.196 2.274 23.500 ;
        RECT 0.000 0.000 1.827 23.500 ;
        LAYER Via1 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal2 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 2.274 0.000 3.167 23.500 ;
        RECT 1.827 0.196 2.274 23.500 ;
        RECT 0.000 0.000 1.827 23.500 ;
        LAYER Via2 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal3 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via3 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal4 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via4 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal5 ;
        RECT 3.467 0.000 4.000 23.500 ;
        RECT 3.167 0.000 3.467 23.350 ;
        RECT 0.000 0.000 3.167 23.500 ;
        LAYER Via5 ;
	RECT 0.000 0.000 4.000 23.500 ;
        LAYER Metal6 ;
        RECT 0.000 0.000 4.000 23.500 ;
    END
END PDO04CDG

MACRO PVDD1DGZ
    CLASS PAD POWER ;
    FOREIGN PVDD1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 23.500 ;
    SYMMETRY x y r90 ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION OUTPUT ;
        USE power ;
        PORT
        LAYER Metal3 ;
        RECT  0.600 22.700 3.400 23.500 ;
        LAYER Metal4 ;
        RECT  0.600 22.700 3.400 23.500 ;
        LAYER Metal5 ;
        RECT  0.600 22.700 3.400 23.500 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 4.000 23.500 ;
#        LAYER Via1 ;
#        RECT  0.5355 22.7480 3.4645 23.2940 ;
#        RECT  2.8820 20.8680 3.4280 22.4540 ;
#        RECT  2.1120 20.8680 2.6580 22.4540 ;
#        RECT  1.3420 20.8680 1.8880 22.4540 ;
#        RECT  0.5720 20.8680 1.1180 22.4540 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 4.000 23.500 ;
#        LAYER Via2 ;
#        RECT  3.4170 23.4570 3.4485 23.4830 ;
#        RECT  0.6165 22.6960 3.4170 23.4830 ;
#        RECT  0.5830 22.6960 0.6165 23.3460 ;
        LAYER Metal3 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
#        LAYER Via3 ;
#        RECT  3.3875 22.7480 3.4645 23.2940 ;
#        RECT  0.5555 22.7480 3.3875 23.4830 ;
#        RECT  0.5355 22.7480 0.5555 23.2940 ;
        LAYER Metal4 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
#        LAYER Via4 ;
#        RECT  3.4170 23.4570 3.4485 23.4830 ;
#        RECT  0.6165 22.6960 3.4170 23.4830 ;
#        RECT  0.5830 22.6960 0.6165 23.3460 ;
        LAYER Metal5 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
#        LAYER Via5 ;
#        RECT  3.3925 22.7430 3.4645 23.2990 ;
#        RECT  0.5505 22.7430 3.3925 23.4880 ;
#        RECT  0.5355 22.7430 0.5505 23.2990 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 4.000 23.500 ;
    END
END PVDD1DGZ

MACRO PVSS1DGZ
    CLASS PAD POWER ;
    FOREIGN PVSS1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 23.500 ;
    SYMMETRY x y r90 ;
    SITE CoreSite ;
    PIN VSS
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
        LAYER Metal3 ;
        RECT  0.600 22.700 3.400 23.500 ;
        LAYER Metal4 ;
        RECT  0.600 22.700 3.400 23.500 ;
        LAYER Metal5 ;
        RECT  0.600 22.700 3.400 23.500 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 4.000 23.500 ;
        LAYER Via1 ;
        RECT  2.8820 20.8680 3.4280 22.4540 ;
        RECT  0.6350 22.7480 3.3650 23.2940 ;
        RECT  2.1120 20.8680 2.6580 22.4540 ;
        RECT  1.3420 20.8680 1.8880 22.4540 ;
        RECT  0.5720 20.8680 1.1180 22.4540 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 4.000 23.500 ;
        LAYER Via2 ;
        RECT  0.6165 23.4570 3.4485 23.4830 ;
        RECT  0.5830 21.8040 3.4170 22.4540 ;
        LAYER Metal3 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
        LAYER Via3 ;
        RECT  0.5555 23.4570 3.3875 23.4830 ;
        LAYER Metal4 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
        LAYER Via4 ;
        RECT  0.6165 23.4570 3.4485 23.4830 ;
        LAYER Metal5 ;
        RECT  3.550 0.000 4.000 23.500 ;
        RECT  0.450 0.000 3.550 22.550 ;
        RECT  0.000 0.000 0.450 23.500 ;
        LAYER Via5 ;
        RECT  0.5505 23.4520 3.3925 23.4880 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 4.000 23.500 ;
    END
END PVSS1DGZ


END LIBRARY

